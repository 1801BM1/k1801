//
// Copyright (c) 2014-2019 by 1801BM1@gmail.com
//______________________________________________________________________________
//
`timescale 1ns / 100ps

module vp_096
(
   input    PIN_CLK,       //
   input    PIN_nINIT,     //
                           //
   input    PIN_nRQ,       //
   input    PIN_nWD,       //
   input    PIN_nCMPC1,    //
   input    PIN_nCMPC2,    //
   input    PIN_nCMPP1,    //
   input    PIN_nCMPP2,    //
                           //
   input    PIN_nDMGIC,    //
   input    PIN_nIAKIC,    //
   output   PIN_nDMGO,     //
   output   PIN_nIAKO,     //
   output   PIN_nDMRC,     //
   output   PIN_nVIRQC,    //
   output   PIN_nSACKC1,   //
   output   PIN_nSACKC2,   //
                           //
   inout    PIN_nSYNCC,    //
   inout    PIN_nDINC,     //
   inout    PIN_nDOUTC,    //
   output   PIN_nWTBTC,    //
   inout    PIN_nRPLYC,    //
   output   PIN_nBSC,      //
                           //
   input    PIN_nSYNCP,    //
   input    PIN_nDINP,     //
   input    PIN_nDOUTP,    //
   input    PIN_nWTBTP,    //
   inout    PIN_nRPLYP,    //
   input    PIN_nBSP,      //
                           //
   output   PIN_CON1,      //
   output   PIN_CON2,      //
   output   PIN_nDLA,      //
   output   PIN_nDLD,      //
   output   PIN_nDLV,      //
   output   PIN_nCLD,      //
   output   PIN_nWWC,      //
   output   PIN_nRDC,      //
   output   PIN_nWWP,      //
   output   PIN_nRDP       //
);

//______________________________________________________________________________
//
// Autogenerated netlist
//
wire CLK2;
wire nSACK_F1;
wire nDMGIC;
wire nSACK_F3;
wire nSACK_F4;
wire SACK_F4;
wire WSELP;
wire WDONE;
wire RDONE;
wire INIT2;
wire nDMGIC_F2;
wire nWD;
wire nDMRC;
wire nCLK2;
wire SACK_F2;
wire nSYNCP1;
wire nINIT;
wire DMRC;
wire RPLYC;
wire WDRQ;
wire INIT1;
wire DLA;
wire nCLD;
wire INIT0;
wire nSYNCC;
wire DOUTP;
wire nIAKIC_F2;
wire nCLK;
wire nWSELC;
wire nSELP;
wire WSELC;
wire DMGIC;
wire nDLV;
wire nSACK_F2;
wire RSELP;
wire SACK_C1;
wire SACK_S1;
wire SACK_F1;
wire BUSYC;
wire nSYNCP0;
wire DINP;
wire INIT3;
wire nIAKIC;
wire IAKIC_F1;
wire DLVD;
wire IRQ;
wire DDONE;
wire CDONE;
wire RSELC;
wire DLD;
wire nVIRQ;
wire VIRQ;
wire nWSELP;
wire nCENA;
wire IAKIC;
wire DINC;
wire SACK_F3;
wire DLV;
wire nSELC;
wire CLK;

wire NET00000, NET00003, NET00007, NET00012, NET00013, NET00014, NET00017, NET00020;
wire NET00021, NET00022, NET00025, NET00026, NET00027, NET00028, NET00029, NET00031;
wire NET00034, NET00035, NET00037, NET00040, NET00041, NET00043, NET00044, NET00045;
wire NET00047, NET00049, NET00051, NET00096, NET00052, NET00054, NET00055, NET00056;
wire NET00057, NET00058, NET00059, NET00061, NET00062, NET00063, NET00064, NET00065;
wire NET00067, NET00068, NET00069, NET00070, NET00072, NET00073, NET00074, NET00076;
wire NET00189, NET00078, NET00079, NET00080, NET00081, NET00082, NET00083, NET00084;
wire NET00085, NET00086, NET00088, NET00090, NET00091, NET00092, NET00093, NET00150;
wire NET00100, NET00101, NET00103, NET00104, NET00105, NET00106, NET00107, NET00110;
wire NET00112, NET00113, NET00114, NET00115, NET00116, NET00117, NET00118, NET00120;
wire NET00121, NET00122, NET00123, NET00124, NET00125, NET00001, NET00127, NET00128;
wire NET00129, NET00130, NET00132, NET00133, NET00135, NET00136, NET00137, NET00138;
wire NET00139, NET00140, NET00141, NET00142, NET00143, NET00144, NET00145, NET00146;
wire NET00147, NET00148, NET00149, NET00152, NET00153, NET00154, NET00157, NET00158;
wire NET00159, NET00160, NET00164, NET00197, NET00198, NET00200, NET00165, NET00201;
wire NET00167, NET00168, NET00169, NET00170, NET00173, NET00175, NET00179, NET00180;
wire NET00181, NET00182, NET00183, NET00184, NET00185, NET00186, NET00187, NET00188;
wire NET00190, NET00191, NET00192, NET00193, NET00194, NET00195, NET00196, NET00202;
wire NET00203, NET00237, NET00239, NET00240, NET00241, NET00243, NET00204, NET00205;
wire NET00206, NET00207, NET00208, NET00209, NET00210, NET00212, NET00213, NET00214;
wire NET00216, NET00217, NET00218, NET00219, NET00221, NET00223, NET00224, NET00225;
wire NET00226, NET00227, NET00228, NET00229, NET00231, NET00232, NET00234, NET00235;
wire NET00263, NET00264, NET00265, NET00266, NET00267, NET00268, NET00292, NET00293;
wire NET00244, NET00245, NET00246, NET00247, NET00248, NET00249, NET00250, NET00251;
wire NET00252, NET00253, NET00254, NET00255, NET00256, NET00257, NET00258, NET00259;
wire NET00260, NET00261, NET00262, NET00294, NET00295, NET00297, NET00301, NET00302;
wire NET00270, NET00269, NET00271, NET00273, NET00274, NET00303, NET00275, NET00276;
wire NET00277, NET00278, NET00279, NET00280, NET00304, NET00282, NET00283, NET00284;
wire NET00285, NET00286, NET00287, NET00288, NET00290, NET00291, NET00305, NET00306;
wire NET00307, NET00309, NET00296, NET00310, NET00298, NET00299, NET00311, NET00308;
wire NET00312;

//______________________________________________________________________________
//
// Autogenerated cell instantiations
//
tOUTPUT_OC cell_PIN15_OC(.x1(NET00055), .y1(PIN_nRPLYC));
tOUTPUT_OC cell_PIN14_OC(.x1(NET00256), .y1(PIN_nSYNCC));
tOUTPUT_OC cell_PIN34_OC(.x1(NET00204), .y1(PIN_nDOUTC));
tOUTPUT_OC cell_PIN3_OC (.x1(nCLD),     .y1(PIN_nDINC));
tOUTPUT_OC cell_PIN23_OC(.x1(NET00190), .y1(PIN_nRPLYP));

tINPUT cell_PIN1 (.y1(NET00054),  .x1(PIN_CLK));
tINPUT cell_PIN41(.y1(NET00041),  .x1(PIN_nINIT));

tOUTPUT cell_PIN11(.x1(NET00049), .y1(PIN_CON2));
tOUTPUT cell_PIN10(.x1(NET00047), .y1(PIN_CON1));
tOUTPUT cell_PIN4 (.x1(nCLD),     .y1(PIN_nCLD));
tOUTPUT cell_PIN8 (.x1(nDLV),     .y1(PIN_nDLV));
tOUTPUT cell_PIN27(.x1(NET00183), .y1(PIN_nDLA));
tOUTPUT cell_PIN29(.x1(NET00192), .y1(PIN_nDLD));
tOUTPUT cell_PIN39(.x1(NET00073), .y1(PIN_nRDP));
tOUTPUT cell_PIN38(.x1(NET00068), .y1(PIN_nRDC));
tOUTPUT cell_PIN40(.x1(NET00133), .y1(PIN_nWWP));
tOUTPUT cell_PIN35(.x1(NET00057), .y1(PIN_nWWC));

tOUTPUT cell_PIN28(.x1(NET00193), .y1(PIN_nWTBTC));
tOUTPUT cell_PIN26(.x1(NET00184), .y1(PIN_nBSC));
tOUTPUT cell_PIN18(.x1(NET00165), .y1(PIN_nDMGO));
tOUTPUT cell_PIN19(.x1(NET00214), .y1(PIN_nSACKC1));
tOUTPUT cell_PIN20(.x1(NET00188), .y1(PIN_nSACKC2));
tOUTPUT cell_PIN7 (.x1(NET00182), .y1(PIN_nIAKO));
tOUTPUT cell_PIN22(.x1(NET00120), .y1(PIN_nDMRC));
tOUTPUT cell_PIN9 (.x1(NET00308), .y1(PIN_nVIRQC));

tINPUT cell_PIN12(.y1(NET00257), .x1(PIN_nDMGIC));
tINPUT cell_PIN15(.y1(NET00248), .x1(PIN_nRPLYC));
tINPUT cell_PIN14(.y1(NET00249), .x1(PIN_nSYNCC));
tINPUT cell_PIN34(.y1(NET00056), .x1(PIN_nDOUTC));
tINPUT cell_PIN2 (.y1(NET00059), .x1(PIN_nIAKIC));
tINPUT cell_PIN3 (.y2(DINC),     .x1(PIN_nDINC));

tINPUT cell_PIN16(.y1(NET00250), .x1(PIN_nSYNCP));
tINPUT cell_PIN25(.y2(NET00179), .x1(PIN_nWTBTP));
tINPUT cell_PIN17(.y2(DOUTP),    .x1(PIN_nDOUTP));
tINPUT cell_PIN24(.y2(NET00180), .x1(PIN_nBSP));
tINPUT cell_PIN5 (.y2(DINP),     .x1(PIN_nDINP));

tINPUT cell_PIN6 (.y1(NET00086), .x1(PIN_nRQ));
tINPUT cell_PIN13(.y1(NET00028), .x1(PIN_nWD));
tINPUT cell_PIN30(.y2(NET00058), .x1(PIN_nCMPC1));
tINPUT cell_PIN31(.y2(NET00061), .x1(PIN_nCMPC2));
tINPUT cell_PIN32(.y2(NET00062), .x1(PIN_nCMPP1));
tINPUT cell_PIN33(.y2(NET00063), .x1(PIN_nCMPP2));

t372 cell_A2(.x1(NET00254), .y2(NET00256), .y3(NET00255), .y4(NET00254), .x5(NET00252), .x6(NET00253));
t372 cell_A14(.x1(NET00144), .y2(NET00146), .y3(NET00145), .y4(NET00144), .x5(RDONE), .x6(NET00146));
t378 cell_A24(.x1(NET00232), .y2(NET00244), .x3(INIT1), .x5(NET00229));
t378 cell_A25(.x1(nCENA), .y2(NET00232), .x3(RDONE), .x5(NET00244));
t379 cell_A29(.x1(NET00246), .y2(NET00247), .x3(INIT2), .y4(NET00245), .x5(NET00245), .x6(nSYNCP1), .x8(NET00247));
t379 cell_A30(.x1(nSYNCP1), .y2(NET00275), .x3(NET00245), .y4(NET00246), .x5(NET00246), .x6(NET00180), .x8(NET00275));
t379 cell_A31(.x1(NET00245), .y2(NET00277), .x3(INIT2), .y4(NET00276), .x5(NET00276), .x6(NET00275), .x8(NET00277));
t379 cell_A35(.x1(NET00278), .y2(NET00283), .x3(INIT2), .y4(NET00279), .x5(NET00279), .x6(nSYNCP1), .x8(NET00283));
t379 cell_A37(.x1(NET00279), .y2(NET00269), .x3(INIT2), .y4(NET00282), .x5(NET00282), .x6(NET00280), .x8(NET00269));
t385 cell_A1(.x1(NET00249), .x2(NET00248), .y3(BUSYC), .x5(NET00248), .y8(RPLYC));
t375 cell_A3(.x1(NET00250), .y2(NET00252), .y3(NET00251), .x4(nSACK_F3), .x5(NET00250), .x6(NET00251), .y9(NET00253));
t378 cell_A26(.x1(NET00229), .y2(NET00228), .x3(RDONE), .x5(NET00232));
t379 cell_A36(.x1(nSYNCP1), .y2(NET00280), .x3(NET00279), .y4(NET00278), .x5(NET00278), .x6(NET00179), .x8(NET00280));
t385 cell_A38(.x1(NET00277), .x2(DLA), .y3(NET00184), .x5(DLA), .y8(NET00183));
t379 cell_C17(.x1(nCLK2), .y2(NET00117), .x3(NET00114), .y4(NET00115), .x5(NET00115), .x6(SACK_F1), .x8(NET00117));
t379 cell_B20(.x1(NET00224), .y2(NET00225), .x3(INIT1), .y4(NET00223), .x5(NET00223), .x6(CLK2), .x8(NET00225));
t375 cell_C20(.x1(NET00213), .y2(NET00214), .y3(NET00118), .x4(SACK_F2), .x5(SACK_F1), .x6(NET00214), .y9(NET00188));
t379 cell_B21(.x1(CLK2), .y2(NET00226), .x3(NET00223), .y4(NET00224), .x5(NET00224), .x6(SACK_F2), .x8(NET00226));
t379 cell_B22(.x1(NET00223), .y2(NET00213), .x3(INIT1), .y4(NET00227), .x5(NET00227), .x6(NET00226), .x8(NET00213));
t378 cell_B25(.x1(NET00231), .y2(CDONE), .x3(NET00232), .x5(INIT1));
t378 cell_B26(.x1(nCENA), .y2(NET00231), .x3(NET00228), .x5(CDONE));
t375 cell_B27(.x1(nCLD), .y2(nCENA), .y3(NET00235), .x4(NET00235), .x5(NET00234), .x6(CDONE), .y9(NET00234));
t372 cell_A16(.x1(NET00147), .y2(NET00149), .y3(NET00148), .y4(NET00147), .x5(NET00145), .x6(NET00149));
t378 cell_B6(.x1(NET00034), .y2(NET00287), .x3(INIT1), .x5(NET00037));
t378 cell_B7(.x1(WDRQ), .y2(NET00034), .x3(DMGIC), .x5(NET00287));
t378 cell_C6(.x1(1'b0), .y2(NET00037), .x3(WDRQ), .x5(NET00035));
t378 cell_C7(.x1(DMRC), .y2(nDMRC), .x3(NET00034), .x5(INIT1));
t378 cell_C8(.x1(WDRQ), .y2(DMRC), .x3(NET00035), .x5(nDMRC));
t378 cell_C11(.x1(1'b0), .y2(NET00113), .x3(SACK_S1), .x5(NET00112));
t378 cell_B11(.x1(NET00110), .y2(NET00138), .x3(INIT1), .x5(NET00113));
t378 cell_B12(.x1(SACK_S1), .y2(NET00110), .x3(SACK_C1), .x5(NET00138));
t378 cell_C12(.x1(nSACK_F1), .y2(SACK_F1), .x3(NET00110), .x5(INIT1));
t391 cell_C14(.x1(nSACK_F1), .x2(NET00118), .y3(NET00312), .y4(NET00120), .x5(nDMRC), .x6(RPLYC), .y9(NET00017), .x10(SACK_F2));
t379 cell_C16(.x1(NET00115), .y2(NET00116), .x3(INIT1), .y4(NET00114), .x5(NET00114), .x6(nCLK2), .x8(NET00116));
t379 cell_C18(.x1(NET00114), .y2(SACK_F2), .x3(INIT1), .y4(NET00121), .x5(NET00121), .x6(NET00117), .x8(SACK_F2));
t378 cell_B24(.x1(1'b0), .y2(NET00229), .x3(nCENA), .x5(NET00228));
t371 cell_J11(.x1(NET00311), .y3(NET00309), .y4(NET00311), .x6(DLVD));
t371 cell_M33(.x1(RSELP), .y3(NET00073), .y4(NET00068), .x6(RSELC));
t378 cell_B8(.x1(NET00037), .y2(NET00035), .x3(DMGIC), .x5(NET00034));
t378 cell_B13(.x1(NET00113), .y2(NET00112), .x3(SACK_C1), .x5(NET00110));
t378 cell_C13(.x1(SACK_S1), .y2(nSACK_F1), .x3(NET00112), .x5(SACK_F1));
t378 cell_C3(.x1(NET00014), .y2(NET00027), .x3(NET00028), .x5(NET00026));
t378 cell_C2(.x1(NET00027), .y2(NET00026), .x3(nSYNCP0), .x5(NET00029));
t428 cell_E6(.x2(INIT0), .y3(INIT1));
t371 cell_D29(.x1(NET00203), .y3(NET00204), .y4(WDONE), .x6(NET00012));
t379 cell_D27(.x1(NET00157), .y2(NET00200), .x3(INIT2), .y4(NET00157), .x5(NET00197), .x6(NET00200), .x8(NET00201));
t383 cell_D8(.x1(NET00312), .y2(SACK_S1), .x3(DMRC), .x4(BUSYC), .x5(nDMGIC), .x6(nDMGIC_F2));
t382 cell_F16(.x1(RDONE), .y2(NET00012), .x3(DDONE), .x4(nSACK_F4), .x5(DOUTP), .x6(NET00013), .y8(NET00013));
t388 cell_F14(.x1(SACK_F4), .y2(RDONE), .x3(nSACK_F2), .y4(DLA), .y5(NET00014), .x6(DMRC), .x7(NET00017), .x10(nINIT));
t379 cell_C4(.x1(nWD), .y2(NET00040), .x3(NET00014), .y4(nWD), .x5(NET00026), .x6(NET00040), .x8(NET00029));
t428 cell_E1(.x2(NET00257), .y3(nDMGIC));
t380 cell_D9(.x1(nDMRC), .y2(NET00165), .y3(NET00164), .x4(nDMGIC_F2), .x5(NET00164), .x6(nDMGIC));
t429 cell_E33(.y3(INIT3), .x5(nINIT));
t428 cell_E8(.x2(NET00121), .y3(nSACK_F2));
t428 cell_K14(.x2(NET00291), .y3(CLK2));
t374 cell_D4(.x1(NET00160), .x2(nDMGIC), .x3(nWD), .y4(WDRQ), .y8(DMGIC));
t378 cell_F3(.x1(nDMGIC), .y2(NET00299), .x3(nDMGIC), .x5(NET00296));
t429 cell_E29(.y3(INIT2), .x5(nINIT));
t379 cell_F24(.x1(NET00150), .y2(NET00152), .x3(INIT2), .y4(NET00150), .x5(nCLK), .x6(NET00152), .x8(NET00153));
t379 cell_C33(.x1(NET00264), .y2(NET00265), .x3(INIT3), .y4(NET00264), .x5(CLK), .x6(NET00265), .x8(NET00266));
t379 cell_F6(.x1(NET00292), .y2(NET00293), .x3(nDMGIC), .y4(NET00292), .x5(nCLK), .x6(NET00293), .x8(NET00294));
t379 cell_F4(.x1(NET00297), .y2(NET00160), .x3(nDMGIC), .y4(NET00297), .x5(NET00296), .x6(NET00160), .x8(NET00298));
t379 cell_F27(.x1(NET00158), .y2(NET00159), .x3(INIT2), .y4(NET00158), .x5(NET00154), .x6(NET00159), .x8(NET00152));
t378 cell_F26(.x1(INIT2), .y2(NET00153), .x3(NET00157), .x5(NET00154));
t378 cell_C35(.x1(INIT3), .y2(NET00266), .x3(NET00158), .x5(NET00267));
t379 cell_C36(.x1(NET00263), .y2(NET00268), .x3(INIT3), .y4(NET00263), .x5(NET00267), .x6(NET00268), .x8(NET00265));
t379 cell_F9(.x1(nDMGIC_F2), .y2(NET00302), .x3(nDMGIC), .y4(nDMGIC_F2), .x5(NET00295), .x6(NET00302), .x8(NET00293));
t378 cell_F8(.x1(nDMGIC), .y2(NET00294), .x3(NET00297), .x5(NET00295));
t379 cell_G38(.x1(nSELP), .y2(NET00243), .x3(INIT3), .y4(nSELP), .x5(NET00241), .x6(NET00243), .x8(NET00239));
t384 cell_F38(.x1(NET00058), .y3(NET00128), .x5(NET00061));
t418 cell_C37(.x1(DLA), .x2(DLD), .y3(NET00192), .y4(NET00193), .x5(NET00269), .x6(NET00179), .x10(DLD));
t379 cell_G9(.x1(NET00043), .y2(DDONE), .x3(nSACK_F2), .y4(NET00051), .x5(NET00051), .x6(NET00052), .x8(DDONE));
t379 cell_D24(.x1(NET00202), .y2(NET00201), .x3(INIT2), .y4(NET00202), .x5(CLK), .x6(NET00201), .x8(NET00198));
t379 cell_F11(.x1(NET00022), .y2(NET00025), .x3(nSACK_F2), .y4(NET00020), .x5(NET00020), .x6(CLK2), .x8(NET00025));
t378 cell_G37(.x1(INIT3), .y2(NET00240), .x3(NET00221), .x5(NET00241));
t378 cell_G36(.x1(NET00240), .y2(NET00241), .x3(nSYNCP1), .x5(NET00239));
t379 cell_F13(.x1(NET00020), .y2(SACK_F3), .x3(nSACK_F2), .y4(nSACK_F3), .x5(nSACK_F3), .x6(NET00021), .x8(SACK_F3));
t378 cell_D26(.x1(INIT2), .y2(NET00198), .x3(WDONE), .x5(NET00197));
t379 cell_C1(.x1(NET00031), .y2(NET00029), .x3(NET00014), .y4(NET00031), .x5(nSYNCP0), .x6(NET00029), .x8(NET00027));
t419 cell_C29(.x1(CDONE), .y2(NET00190), .x4(NET00136), .x5(NET00148), .x6(DOUTP), .x10(DDONE));
t387 cell_D34(.x1(NET00263), .y2(DLD), .x3(NET00158), .y4(NET00203), .x5(NET00158), .x6(NET00263));
t379 cell_F1(.x1(NET00301), .y2(NET00298), .x3(nDMGIC), .y4(NET00301), .x5(CLK), .x6(NET00298), .x8(NET00299));
t382 cell_D11(.x1(BUSYC), .y2(NET00096), .x3(DMGIC), .x4(nDMRC), .x5(NET00096), .x6(nSACK_F4), .y8(SACK_C1));
t428 cell_K13(.x2(NET00290), .y3(nCLK2));
t428 cell_K22(.x2(NET00041), .y3(nINIT));
t378 cell_F25(.x1(NET00153), .y2(NET00154), .x3(nCLK), .x5(NET00152));
t378 cell_C34(.x1(NET00266), .y2(NET00267), .x3(CLK), .x5(NET00265));
t378 cell_F7(.x1(NET00294), .y2(NET00295), .x3(nCLK), .x5(NET00293));
t379 cell_F12(.x1(CLK2), .y2(NET00021), .x3(NET00020), .y4(NET00022), .x5(NET00022), .x6(SACK_F2), .x8(NET00021));
t378 cell_D25(.x1(NET00198), .y2(NET00197), .x3(CLK), .x5(NET00201));
t379 cell_G35(.x1(NET00237), .y2(NET00239), .x3(INIT3), .y4(NET00237), .x5(nSYNCP1), .x6(NET00239), .x8(NET00240));
t379 cell_G7(.x1(NET00044), .y2(NET00045), .x3(nSACK_F2), .y4(NET00043), .x5(NET00043), .x6(DLD), .x8(NET00045));
t379 cell_G8(.x1(DLD), .y2(NET00052), .x3(NET00043), .y4(NET00044), .x5(NET00044), .x6(1'b1), .x8(NET00052));
t389 cell_I30(.x1(NET00208), .x2(RSELC), .y3(NET00055), .x4(NET00209), .y5(NET00057), .x6(NET00194), .x10(NET00092));
t379 cell_I33(.x1(NET00206), .y2(NET00207), .x3(nWSELP), .y4(NET00205), .x5(NET00205), .x6(CLK2), .x8(NET00207));
t379 cell_I35(.x1(NET00205), .y2(NET00106), .x3(nWSELP), .y4(NET00212), .x5(NET00212), .x6(NET00210), .x8(NET00106));
t379 cell_J29(.x1(NET00065), .y2(NET00067), .x3(nWSELC), .y4(NET00064), .x5(NET00064), .x6(CLK2), .x8(NET00067));
t380 cell_L4(.x1(DINC), .y2(IAKIC), .y3(NET00170), .x4(VIRQ), .x5(nIAKIC), .x6(IAKIC));
t386 cell_J4(.x1(nDLV), .y2(NET00307), .y3(DLVD), .y4(NET00308), .x5(VIRQ), .x6(DLV), .x7(NET00307));
t382 cell_L8(.x1(nIAKIC_F2), .y2(NET00173), .x3(nVIRQ), .x4(nIAKIC), .x5(NET00170), .x6(DLVD), .y8(NET00175));
t372 cell_B1(.x1(NET00249), .y2(NET00167), .y3(NET00286), .y4(NET00285), .x5(NET00285), .x6(NET00286));
t379 cell_L34(.x1(CLK2), .y2(NET00141), .x3(NET00140), .y4(NET00142), .x5(NET00142), .x6(NET00103), .x8(NET00141));
t379 cell_L33(.x1(NET00142), .y2(NET00143), .x3(nWSELP), .y4(NET00140), .x5(NET00140), .x6(CLK2), .x8(NET00143));
t379 cell_J24(.x1(NET00083), .y2(NET00084), .x3(nWSELC), .y4(NET00082), .x5(NET00082), .x6(nCLK2), .x8(NET00084));
t378 cell_L1(.x1(NET00186), .y2(NET00187), .x3(INIT0), .x5(NET00185));
t378 cell_M8(.x1(nIAKIC), .y2(NET00261), .x3(NET00070), .x5(NET00258));
t379 cell_H13(.x1(NET00000), .y2(SACK_F4), .x3(nSACK_F2), .y4(nSACK_F4), .x5(nSACK_F4), .x6(NET00007), .x8(SACK_F4));
t379 cell_H12(.x1(nCLK2), .y2(NET00007), .x3(NET00000), .y4(NET00001), .x5(NET00001), .x6(SACK_F3), .x8(NET00007));
t379 cell_N33(.x1(NET00105), .y2(NET00107), .x3(nWSELP), .y4(NET00101), .x5(NET00101), .x6(nCLK2), .x8(NET00107));
t388 cell_M34(.x1(RSELP), .y2(NET00136), .x3(NET00135), .y4(NET00137), .y5(NET00133), .x6(NET00106), .x7(NET00137), .x10(NET00100));
t379 cell_L35(.x1(NET00140), .y2(NET00135), .x3(nWSELP), .y4(NET00139), .x5(NET00139), .x6(NET00141), .x8(NET00135));
t379 cell_J26(.x1(NET00082), .y2(NET00092), .x3(nWSELC), .y4(NET00091), .x5(NET00091), .x6(NET00088), .x8(NET00092));
t378 cell_L3(.x1(NET00185), .y2(NET00191), .x3(IAKIC), .x5(NET00186));
t378 cell_M1(.x1(1'b0), .y2(NET00185), .x3(NET00189), .x5(NET00191));
t378 cell_M7(.x1(NET00261), .y2(NET00258), .x3(nCLK), .x5(NET00260));
t428 cell_K11(.x2(NET00054), .y3(CLK));
t379 cell_H24(.x1(NET00132), .y2(NET00130), .x3(INIT3), .y4(NET00132), .x5(nSYNCC), .x6(NET00130), .x8(NET00127));
t378 cell_H25(.x1(NET00127), .y2(NET00125), .x3(nSYNCC), .x5(NET00130));
t428 cell_K6(.x2(NET00059), .y3(nIAKIC));
t429 cell_K24(.y3(INIT0), .x5(NET00041));
t379 cell_N35(.x1(NET00101), .y2(NET00103), .x3(nWSELP), .y4(NET00100), .x5(NET00100), .x6(NET00104), .x8(NET00103));
t378 cell_M3(.x1(NET00189), .y2(nVIRQ), .x3(NET00191), .x5(VIRQ));
t378 cell_M2(.x1(nVIRQ), .y2(VIRQ), .x3(NET00186), .x5(INIT0));
t377 cell_J27(.x1(NET00093), .y2(nWSELC), .x3(nSELC), .y4(RSELC), .x5(WSELC), .x6(NET00056), .x8(nSELC), .y9(WSELC));
t372 cell_J12(.x1(DINC), .y2(NET00310), .y3(NET00093), .y4(NET00208), .x5(NET00309), .x6(NET00310));
t379 cell_H29(.x1(NET00123), .y2(NET00124), .x3(nWSELC), .y4(NET00122), .x5(NET00122), .x6(nCLK2), .x8(NET00124));
t379 cell_H27(.x1(nSELC), .y2(NET00129), .x3(INIT3), .y4(nSELC), .x5(NET00125), .x6(NET00129), .x8(NET00130));
t429 cell_K9(.y3(nCLK), .x5(NET00054));
t387 cell_N2(.x1(nINIT), .y2(NET00079), .x3(IRQ), .y4(NET00189), .x5(nVIRQ), .x6(IAKIC_F1));
t372 cell_H6(.x1(NET00168), .y2(NET00169), .y3(nSYNCC), .y4(NET00168), .x5(NET00167), .x6(NET00169));
t379 cell_J9(.x1(NET00290), .y2(NET00291), .x3(INIT0), .y4(NET00290), .x5(NET00303), .x6(NET00291), .x8(NET00305));
t379 cell_O6(.x1(NET00076), .y2(NET00072), .x3(nIAKIC), .y4(NET00076), .x5(CLK), .x6(NET00072), .x8(NET00074));
t378 cell_L13(.x1(NET00271), .y2(NET00270), .x3(NET00175), .x5(NET00273));
t378 cell_O7(.x1(NET00074), .y2(NET00069), .x3(CLK), .x5(NET00072));
t378 cell_L12(.x1(NET00173), .y2(NET00273), .x3(NET00175), .x5(NET00274));
t379 cell_H31(.x1(NET00122), .y2(NET00209), .x3(nWSELC), .y4(NET00216), .x5(NET00216), .x6(NET00217), .x8(NET00209));
t379 cell_H30(.x1(nCLK2), .y2(NET00217), .x3(NET00122), .y4(NET00123), .x5(NET00123), .x6(NET00195), .x8(NET00217));
t384 cell_I6(.x1(DINP), .y3(nCLD), .x5(SACK_F4));
t379 cell_O9(.x1(NET00070), .y2(IAKIC_F1), .x3(nIAKIC), .y4(NET00070), .x5(NET00069), .x6(IAKIC_F1), .x8(NET00072));
t379 cell_O3(.x1(NET00078), .y2(NET00080), .x3(NET00079), .y4(IRQ), .x5(IRQ), .x6(NET00081), .x8(NET00080));
t378 cell_O8(.x1(nIAKIC), .y2(NET00074), .x3(nIAKIC), .x5(NET00069));
t378 cell_M11(.x1(1'b0), .y2(NET00271), .x3(NET00173), .x5(NET00270));
t378 cell_M12(.x1(nDLV), .y2(DLV), .x3(NET00273), .x5(INIT0));
t386 cell_H35(.x1(NET00062), .y2(NET00219), .y3(NET00218), .y4(NET00221), .x5(NET00063), .x6(DINP), .x7(DOUTP));
t378 cell_J8(.x1(INIT0), .y2(NET00304), .x3(NET00291), .x5(NET00303));
t379 cell_O1(.x1(NET00085), .y2(NET00090), .x3(NET00079), .y4(NET00078), .x5(NET00078), .x6(NET00086), .x8(NET00090));
t379 cell_O2(.x1(NET00086), .y2(NET00081), .x3(NET00078), .y4(NET00085), .x5(NET00085), .x6(1'b1), .x8(NET00081));
t378 cell_F2(.x1(NET00299), .y2(NET00296), .x3(CLK), .x5(NET00298));
t382 cell_G6(.x1(DLV), .y2(NET00047), .x3(DLA), .x4(RSELC), .x5(NET00047), .x6(DLD), .y8(NET00049));
t379 cell_H11(.x1(NET00001), .y2(NET00003), .x3(nSACK_F2), .y4(NET00000), .x5(NET00000), .x6(nCLK2), .x8(NET00003));
t379 cell_I34(.x1(CLK2), .y2(NET00210), .x3(NET00205), .y4(NET00206), .x5(NET00206), .x6(WSELP), .x8(NET00210));
t379 cell_N34(.x1(nCLK2), .y2(NET00104), .x3(NET00101), .y4(NET00105), .x5(NET00105), .x6(NET00106), .x8(NET00104));
t379 cell_J30(.x1(CLK2), .y2(NET00196), .x3(NET00064), .y4(NET00065), .x5(NET00065), .x6(NET00092), .x8(NET00196));
t379 cell_J25(.x1(nCLK2), .y2(NET00088), .x3(NET00082), .y4(NET00083), .x5(NET00083), .x6(WSELC), .x8(NET00088));
t380 cell_L6(.x1(nIAKIC_F2), .y2(NET00182), .y3(NET00181), .x4(nIAKIC), .x5(NET00181), .x6(VIRQ));
t379 cell_J6(.x1(NET00306), .y2(NET00305), .x3(INIT0), .y4(NET00306), .x5(CLK), .x6(NET00305), .x8(NET00304));
t378 cell_L2(.x1(NET00189), .y2(NET00186), .x3(IAKIC), .x5(NET00187));
t377 cell_H34(.x1(NET00218), .y2(nWSELP), .x3(nSELP), .y4(WSELP), .x5(WSELP), .x6(nSELP), .x8(NET00219), .y9(RSELP));
t378 cell_H26(.x1(INIT3), .y2(NET00127), .x3(NET00128), .x5(NET00125));
t379 cell_J31(.x1(NET00064), .y2(NET00195), .x3(nWSELC), .y4(NET00194), .x5(NET00194), .x6(NET00196), .x8(NET00195));
t379 cell_M9(.x1(nIAKIC_F2), .y2(NET00259), .x3(nIAKIC), .y4(nIAKIC_F2), .x5(NET00258), .x6(NET00259), .x8(NET00260));
t378 cell_J7(.x1(NET00304), .y2(NET00303), .x3(CLK), .x5(NET00305));
t379 cell_M6(.x1(NET00262), .y2(NET00260), .x3(nIAKIC), .y4(NET00262), .x5(nCLK), .x6(NET00260), .x8(NET00261));
t378 cell_M13(.x1(NET00173), .y2(nDLV), .x3(NET00270), .x5(DLV));
t378 cell_L11(.x1(NET00273), .y2(NET00274), .x3(INIT0), .x5(NET00271));
t371 cell_B2(.x1(NET00255), .y3(NET00284), .y4(nSYNCP0), .x6(NET00284));
t371 cell_B4(.x1(NET00288), .y3(nSYNCP1), .y4(NET00288), .x6(NET00255));

endmodule
