//
// Copyright (c) 2013-2014 by 1801BM1@gmail.com
//______________________________________________________________________________
//
`timescale 1ns / 100ps

module vp_014
(
   inout[7:0]  PIN_nAD,       // Address/Data inverted bus
                              //
   input       PIN_nSYNC,     //
   input       PIN_nDIN,      //
   input       PIN_nDOUT,     //
   input       PIN_nINIT,     //
   input       PIN_nCS,       //
   input       PIN_nIAKI,     //
   output      PIN_nIAKO,     //
   output      PIN_nRPLY,     //
   output      PIN_nIRQ,      //
                              //
   input[7:1]  PIN_Y,         //
   output[7:1] PIN_Y_OC,      //
   input[9:0]  PIN_X,         //
   output      PIN_RP1_OC,    //
   output      PIN_RP2_OC,    //
   input       PIN_RP1,       //
   input       PIN_RP2,       //
                              //
   input       PIN_nCTRL,     //
   input       PIN_nSHIFT,    //
   input       PIN_nEC1,      //
   input       PIN_EC2        //
);

//______________________________________________________________________________
//
// Autogenerated netlist
//
wire nSYNC;
wire nCTRL;

wire nC0;
wire nC1;
wire nC2;
wire nC3;
wire nC4;
wire C5;
wire C6;

wire X0;
wire X1;
wire X2;
wire X3;
wire X4;
wire X5;
wire X6;
wire X7;
wire X8;
wire X9;
wire nX5;
wire nX4X5;

wire Y1IN;
wire Y3IN;
wire Y4IN;
wire Y5IN;
wire Y6IN;
wire Y7IN;
wire Y2IN;

wire nY1OC;
wire nY2OC;
wire nY3OC;
wire nY5OC;

wire nX6_9;
wire X0_3;

wire nV274;
wire nLOCK;
wire RP2;
wire XANY;
wire nREADY;
wire LOCK;
wire RELEASE;
wire WSTB;
wire SHIFT;
wire IEN;
wire nDIN;
wire DATRD;
wire IACK;
wire VANY;
wire nOE;
wire nCSR;
wire nEC2;
wire EC1;
wire nIEN;
wire nIRQ;
wire INIT;
wire nXANY;
wire READY;
wire nCSRRD;
wire PRESS;
wire BUSY;
wire nCSRWR;
wire nDAT;

wire NET00225;
wire NET00006;
wire NET00008;
wire NET00010;
wire NET00013;
wire NET00014;
wire NET00015;
wire NET00016;
wire NET00017;
wire NET00018;
wire NET00021;
wire NET00022;
wire NET00023;
wire NET00024;
wire NET00183;
wire NET00026;
wire NET00028;
wire NET00090;
wire NET00031;
wire NET00188;
wire NET00034;
wire NET00186;
wire NET00037;
wire NET00187;
wire NET00039;
wire NET00121;
wire NET00041;
wire NET00042;
wire NET00100;
wire NET00046;
wire NET00047;
wire NET00109;
wire NET00050;
wire NET00052;
wire NET00053;
wire NET00058;
wire NET00060;
wire NET00061;
wire NET00062;
wire NET00063;
wire NET00064;
wire NET00065;
wire NET00066;
wire NET00067;
wire NET00068;
wire NET00069;
wire NET00070;
wire NET00072;
wire NET00002;
wire NET00076;
wire NET00077;
wire NET00079;
wire NET00080;
wire NET00082;
wire NET00084;
wire NET00087;
wire NET00088;
wire NET00089;
wire NET00101;
wire NET00092;
wire NET00095;
wire NET00098;
wire NET00099;
wire NET00106;
wire NET00193;
wire NET00102;
wire NET00104;
wire NET00105;
wire NET00181;
wire NET00107;
wire NET00108;
wire NET00210;
wire NET00110;
wire NET00223;
wire NET00113;
wire NET00114;
wire NET00117;
wire NET00118;
wire NET00119;
wire NET00209;
wire NET00122;
wire NET00123;
wire NET00124;
wire NET00128;
wire NET00130;
wire NET00132;
wire NET00133;
wire NET00135;
wire NET00136;
wire NET00137;
wire NET00139;
wire NET00140;
wire NET00197;
wire NET00145;
wire NET00205;
wire NET00147;
wire NET00204;
wire NET00151;
wire NET00152;
wire NET00153;
wire NET00154;
wire NET00155;
wire NET00156;
wire NET00158;
wire NET00159;
wire NET00191;
wire NET00164;
wire NET00166;
wire NET00167;
wire NET00168;
wire NET00169;
wire NET00170;
wire NET00171;
wire NET00172;
wire NET00173;
wire NET00174;
wire NET00175;
wire NET00176;
wire NET00177;
wire NET00178;
wire NET00179;
wire NET00195;
wire NET00182;
wire NET00184;
wire NET00185;
wire NET00198;
wire NET00206;
wire NET00196;
wire NET00203;
wire NET00211;
wire NET00215;
wire NET00194;
wire NET00214;
wire NET00222;
wire NET00221;
wire NET00212;
wire NET00199;
wire NET00200;
wire NET00201;
wire NET00202;
wire NET00213;
wire NET00217;
wire NET00218;
wire NET00220;
wire NET00219;

//______________________________________________________________________________
//
// Autogenerated cell instantiations
//
tOUTPUT_OE cell_PINOU39(.x1(NET00107), .x2(NET00076), .y1(PIN_nAD[0]));
tOUTPUT_OE cell_PINOU32(.x1(NET00110), .x2(NET00076), .y1(PIN_nAD[1]));
tOUTPUT_OE cell_PINOU37(.x1(NET00102), .x2(NET00076), .y1(PIN_nAD[2]));
tOUTPUT_OE cell_PINOU36(.x1(NET00223), .x2(NET00076), .y1(PIN_nAD[3]));
tOUTPUT_OE cell_PINOU35(.x1(NET00185), .x2(NET00076), .y1(PIN_nAD[4]));
tOUTPUT_OE cell_PINOU34(.x1(NET00183), .x2(NET00076), .y1(PIN_nAD[5]));
tOUTPUT_OE cell_PINOU33(.x1(NET00090), .x2(NET00076), .y1(PIN_nAD[6]));
tOUTPUT_OE cell_PINOU38(.x1(NET00188), .x2(NET00076), .y1(PIN_nAD[7]));

tINPUT cell_PIN32(.y1(NET00079), .x1(PIN_nAD[1]));
tINPUT cell_PIN33(.y1(NET00080), .x1(PIN_nAD[6]));

tINPUT cell_PIN15(.y2(X0), .x1(PIN_X[0]));
tINPUT cell_PIN14(.y2(X1), .x1(PIN_X[1]));
tINPUT cell_PIN13(.y2(X2), .x1(PIN_X[2]));
tINPUT cell_PIN12(.y2(X3), .x1(PIN_X[3]));
tINPUT cell_PIN11(.y2(X4), .x1(PIN_X[4]));
tINPUT cell_PIN10(.y2(X5), .x1(PIN_X[5]));
tINPUT cell_PIN9( .y2(X6), .x1(PIN_X[6]));
tINPUT cell_PIN8( .y2(X7), .x1(PIN_X[7]));
tINPUT cell_PIN7( .y2(X8), .x1(PIN_X[8]));
tINPUT cell_PIN6( .y2(X9), .x1(PIN_X[9]));

tINPUT cell_PIN5( .y2(NET00193), .x1(PIN_Y[1]));
tINPUT cell_PIN4( .y2(NET00028), .x1(PIN_Y[2]));
tINPUT cell_PIN3( .y2(NET00181), .x1(PIN_Y[3]));
tINPUT cell_PIN2( .y2(NET00210), .x1(PIN_Y[4]));
tINPUT cell_PIN1( .y2(NET00209), .x1(PIN_Y[5]));
tINPUT cell_PIN41(.y2(NET00026), .x1(PIN_Y[6]));
tINPUT cell_PIN40(.y2(NET00023), .x1(PIN_Y[7]));

tOUTPUT cell_PIN24(.x1(NET00167), .y1(PIN_nIAKO));

tOUTPUT_OC cell_PIN5_OC( .x1(nY1OC),   .y1(PIN_Y_OC[1]));
tOUTPUT_OC cell_PIN4_OC( .x1(nY2OC),   .y1(PIN_Y_OC[2]));
tOUTPUT_OC cell_PIN3_OC( .x1(nY3OC),   .y1(PIN_Y_OC[3]));
tOUTPUT_OC cell_PIN2_OC( .x1(NET00203),.y1(PIN_Y_OC[4]));
tOUTPUT_OC cell_PIN1_OC( .x1(nY5OC),   .y1(PIN_Y_OC[5]));
tOUTPUT_OC cell_PIN41_OC(.x1(NET00024),.y1(PIN_Y_OC[6]));
tOUTPUT_OC cell_PIN40_OC(.x1(NET00022),.y1(PIN_Y_OC[7]));

tOUTPUT_OC cell_PIN23_OC(.x1(NET00225),.y1(PIN_nIRQ));
tOUTPUT_OC cell_PIN28_OC(.x1(NET00196),.y1(PIN_nRPLY));
tOUTPUT_OC cell_PIN20_OC(.x1(XANY),    .y1(PIN_RP1_OC));
tOUTPUT_OC cell_PIN22_OC(.x1(nXANY),   .y1(PIN_RP2_OC));

tINPUT cell_PIN16(.y1(SHIFT),    .x1(PIN_nSHIFT));
tINPUT cell_PIN17(.y1(EC1),      .x1(PIN_nEC1));
tINPUT cell_PIN31(.y2(nEC2),     .x1(PIN_EC2));
tINPUT cell_PIN18(.y2(nCTRL),    .x1(PIN_nCTRL));
tINPUT cell_PIN19(.y2(INIT),     .x1(PIN_nINIT));
tINPUT cell_PIN25(.y1(NET00124), .x1(PIN_nIAKI));
tINPUT cell_PIN29(.y1(NET00171), .x1(PIN_nSYNC));
tINPUT cell_PIN27(.y1(NET00168), .x1(PIN_nDOUT));
tINPUT cell_PIN30(.y2(NET00077), .x1(PIN_nCS));
tINPUT cell_PIN26(.y1(nDIN),     .x1(PIN_nDIN));
tINPUT cell_PIN20(.y2(NET00170), .x1(PIN_RP1));
tINPUT cell_PIN22(.y2(NET00058), .x1(PIN_RP2));

//______________________________________________________________________________
//
t370 cell_I33(.y2(NET00179), .x5(NET00168));
t428 cell_E31(.x2(LOCK), .y3(NET00021));
t428 cell_E33(.x2(NET00171), .y3(nSYNC));
t373 cell_I7(.x1(NET00201), .x3(DATRD), .y4(NET00199));
t379 cell_H7(.x1(READY), .y2(NET00159), .x3(INIT), .y4(BUSY), .x5(BUSY), .x6(RELEASE), .x8(NET00159));
t429 cell_E3(.y3(NET00101), .x5(DATRD));
t381 cell_H17(.x1(X9), .y2(nC3), .x3(NET00013), .x4(NET00015), .x6(NET00014));
t381 cell_H18(.x1(Y4IN), .y2(nC2), .x3(Y5IN), .x4(Y7IN), .x6(Y6IN));
t416 cell_D33(.c1(nSYNC), .q3(NET00204), .q4(NET00205), .d5(NET00079));
t382 cell_F29(.x1(NET00152), .y2(NET00154), .x3(NET00153), .x4(NET00155), .x5(NET00151), .x6(X0), .y8(NET00152));
t371 cell_G0(.x1(NET00070), .y3(NET00063), .y4(NET00070), .x6(NET00068));
t382 cell_C11(.x1(DATRD), .y2(nOE), .x3(NET00117), .x4(NET00113), .x5(nV274), .x6(NET00118), .y8(NET00118));
t371 cell_F1(.x1(NET00220), .y3(NET00069), .y4(NET00220), .x6(NET00219));
t388 cell_L15(.x1(nX4X5), .y2(NET00214), .x3(NET00213), .y4(NET00017), .y5(NET00212), .x6(SHIFT), .x7(NET00047), .x10(NET00214));
t391 cell_F31(.x1(X2), .x2(NET00197), .y3(NET00153), .y4(NET00197), .x5(Y1IN), .x6(Y1IN), .y9(NET00151), .x10(X1));
t384 cell_F33(.x1(NET00179), .y3(nCSRWR), .x5(NET00198));
t428 cell_E11(.x2(nOE), .y3(NET00076));
t379 cell_D11(.x1(NET00092), .y2(IEN), .x3(INIT), .y4(nIEN), .x5(nIEN), .x6(NET00095), .x8(IEN));
t379 cell_G3(.x1(NET00061), .y2(NET00066), .x3(NET00062), .y4(NET00061), .x5(RP2), .x6(NET00066), .x8(NET00063));
t371 cell_G1(.x1(NET00067), .y3(NET00068), .y4(NET00067), .x6(NET00069));
t378 cell_C18(.x1(NET00124), .y2(IACK), .x3(nDIN), .x5(NET00123));
t379 cell_I17(.x1(X8), .y2(NET00015), .x3(X6), .y4(NET00014), .x5(nX5), .x6(NET00006), .x8(X8));
t374 cell_G27(.x1(NET00132), .x2(nX4X5), .x3(NET00139), .y4(NET00140), .y8(NET00139));
t377 cell_H26(.x1(nCTRL), .y2(NET00130), .x3(NET00130), .y4(NET00132), .x5(NET00128), .x6(SHIFT), .x8(nX6_9), .y9(NET00133));
t374 cell_G9(.x1(PRESS), .x2(RP2), .x3(NET00072), .y4(RELEASE), .y8(NET00065));
t373 cell_J5(.x1(BUSY), .x3(RELEASE), .y4(NET00200));
t379 cell_I5(.x1(NET00200), .y2(NET00202), .x3(INIT), .y4(NET00201), .x5(NET00201), .x6(DATRD), .x8(NET00202));
t370 cell_F11(.y2(nX5), .x5(X5));
t381 cell_I18(.x1(X8), .y2(NET00013), .x3(X6), .x4(NET00037), .x6(X4));
t378 cell_L17(.x1(nY3OC), .y2(NET00215), .x3(Y4IN), .x5(Y5IN));
t416 cell_H33(.c1(nSYNC), .q4(NET00191), .d5(NET00077));
t391 cell_G30(.x1(X0), .x2(NET00194), .y3(NET00155), .y4(NET00175), .x5(Y3IN), .x6(Y3IN), .y9(NET00194), .x10(X1));
t371 cell_C7(.x1(nXANY), .y3(XANY), .y4(RP2), .x6(NET00058));
t379 cell_I9(.x1(nREADY), .y2(READY), .x3(NET00199), .y4(nREADY), .x5(INIT), .x6(READY), .x8(NET00200));
t376 cell_L5(.x1(NET00164), .x3(nREADY), .y4(NET00166), .x6(IACK), .x8(NET00166), .y9(NET00164));
t390 cell_M17(.x1(NET00203), .y4(Y4IN), .x5(NET00210), .x6(NET00021), .y9(NET00203), .x10(Y4IN));
t390 cell_M19(.x1(nY5OC), .y4(Y5IN), .x5(NET00209), .x6(NET00021), .y9(nY5OC), .x10(Y5IN));
t390 cell_H31(.x1(nY1OC), .y4(Y1IN), .x5(NET00193), .x6(NET00021), .y9(nY1OC), .x10(Y1IN));
t373 cell_I11(.x1(X5), .x3(X4), .y4(nX4X5));
t376 cell_D9(.x1(NET00080), .x3(nCSRWR), .y4(NET00092), .x6(nCSRWR), .x8(NET00092), .y9(NET00095));
t370 cell_H11(.y2(NET00006), .x5(X7));
t373 cell_F20(.x1(nLOCK), .x3(INIT), .y4(LOCK));
t376 cell_C21(.x1(NET00034), .x3(NET00101), .y4(NET00182), .x6(VANY), .x8(NET00182), .y9(NET00183));
t381 cell_J21(.x1(nY1OC), .y2(NET00082), .x3(Y2IN), .x4(Y6IN), .x6(Y4IN));
t379 cell_L21(.x1(Y6IN), .y2(NET00050), .x3(Y4IN), .y4(NET00052), .x5(nY3OC), .x6(Y6IN), .x8(nY5OC));
t370 cell_D13(.y2(NET00087), .x5(X4));
t379 cell_G7(.x1(NET00062), .y2(NET00064), .x3(NET00063), .y4(NET00062), .x5(NET00061), .x6(NET00064), .x8(NET00065));
t379 cell_F9(.x1(PRESS), .y2(NET00156), .x3(NET00061), .y4(PRESS), .x5(RP2), .x6(NET00156), .x8(NET00064));
t387 cell_L11(.x1(nX4X5), .y2(NET00217), .x3(NET00217), .y4(nXANY), .x5(nX6_9), .x6(X0_3));
t416 cell_F23(.c1(NET00145), .q3(NET00122), .d5(NET00002));
t381 cell_I23(.x1(X9), .y2(NET00018), .x3(NET00084), .x4(NET00088), .x6(X8));
t374 cell_I24(.x1(NET00101), .x2(NET00108), .x3(NET00109), .y4(NET00108), .y8(NET00110));
t381 cell_F13(.x1(X3), .y2(NET00053), .x3(X1), .x4(X2), .x6(X0));
t373 cell_G13(.x1(X3), .x3(X1), .y4(NET00037));
t416 cell_C23(.c1(nDIN), .q3(NET00123), .q4(NET00178), .d5(NET00060));
t374 cell_D23(.x1(NET00154), .x2(NET00175), .x3(NET00176), .y4(NET00174), .y8(NET00176));
t374 cell_I25(.x1(NET00101), .x2(NET00105), .x3(NET00106), .y4(NET00105), .y8(NET00107));
t381 cell_I26(.x1(X9), .y2(NET00104), .x3(X7), .x4(X6), .x6(X8));
t391 cell_J13(.x1(NET00212), .x2(SHIFT), .y3(NET00222), .y4(NET00213), .x5(NET00221), .x6(NET00047), .y9(NET00221), .x10(NET00222));
t377 cell_C29(.x1(NET00186), .y2(NET00186), .x3(NET00187), .y4(NET00188), .x5(nV274), .x6(nREADY), .x8(nCSRRD), .y9(NET00187));
t390 cell_I30(.x1(nY3OC), .y4(Y3IN), .x5(NET00181), .x6(NET00021), .y9(nY3OC), .x10(Y3IN));
t376 cell_C25(.x1(NET00101), .x3(NET00039), .y4(NET00184), .x6(NET00184), .x8(VANY), .y9(NET00185));
t428 cell_E17(.x2(WSTB), .y3(NET00145));
t390 cell_C33(.x1(NET00204), .y4(nDAT), .x5(NET00191), .x6(NET00205), .y9(nCSR), .x10(NET00191));
t373 cell_D25(.x1(nEC2), .x3(NET00174), .y4(NET00002));
t378 cell_J25(.x1(NET00087), .y2(NET00088), .x3(X6), .x5(X7));
t381 cell_L23(.x1(Y4IN), .y2(NET00046), .x3(Y5IN), .x4(Y7IN), .x6(Y6IN));
t416 cell_G16(.c1(NET00145), .q3(NET00031), .d5(C6));
t373 cell_G25(.x1(NET00104), .x3(nCTRL), .y4(C6));
t380 cell_G23(.x1(NET00140), .y2(X0_3), .y3(C5), .x4(NET00133), .x5(NET00053), .x6(X0_3));
t390 cell_M25(.x1(NET00024), .y4(Y6IN), .x5(NET00026), .x6(NET00021), .y9(NET00024), .x10(Y6IN));
t390 cell_M23(.x1(nY2OC), .y4(Y2IN), .x5(NET00028), .x6(NET00021), .y9(nY2OC), .x10(Y2IN));
t416 cell_G19(.c1(NET00145), .q4(NET00041), .d5(nC3));
t381 cell_H21(.x1(NET00050), .y2(nC0), .x3(NET00052), .x4(Y7IN), .x6(NET00082));
t373 cell_L25(.x1(nX5), .x3(NET00046), .y4(NET00047));
t416 cell_G21(.c1(NET00145), .q4(NET00109), .d5(nC1));
t380 cell_D31(.x1(nDIN), .y2(NET00206), .y3(DATRD), .x4(nDAT), .x5(nDIN), .x6(nSYNC));
t385 cell_L31(.x1(NET00147), .x2(EC1), .y3(NET00136), .x5(NET00042), .y8(NET00147));
t376 cell_H16(.x1(NET00010), .x3(NET00016), .y4(nC4), .x6(NET00017), .x8(NET00018), .y9(NET00016));
t391 cell_M31(.x1(NET00135), .x2(NET00042), .y3(NET00135), .y4(NET00137), .x5(EC1), .x6(NET00137), .y9(NET00128), .x10(NET00136));
t370 cell_H23(.y2(NET00098), .x5(nV274));
t376 cell_H9(.x1(PRESS), .x3(NET00158), .y4(NET00072), .x6(NET00159), .x8(NET00072), .y9(NET00158));
t373 cell_H5(.x1(nIEN), .x3(nIRQ), .y4(NET00060));
t374 cell_C13(.x1(IEN), .x2(nCSRRD), .x3(nCSRRD), .y4(NET00114), .y8(NET00113));
t374 cell_L7(.x1(nREADY), .x2(NET00169), .x3(NET00166), .y4(NET00169), .y8(nIRQ));
t371 cell_F0(.x1(NET00218), .y3(NET00219), .y4(NET00218), .x6(NET00170));
t381 cell_H19(.x1(NET00211), .y2(nC1), .x3(NET00215), .x4(Y7IN), .x6(Y6IN));
t385 cell_C17(.x1(nV274), .x2(NET00119), .y3(VANY), .x5(NET00119), .y8(NET00117));
t378 cell_L19(.x1(Y5IN), .y2(NET00211), .x3(Y4IN), .x5(nY2OC));
t385 cell_G33(.x1(nCSRWR), .x2(NET00195), .y3(NET00195), .x5(NET00076), .y8(NET00196));
t370 cell_C9(.y2(NET00225), .x5(NET00060));
t376 cell_D7(.x1(PRESS), .x3(XANY), .y4(nLOCK), .x6(NET00156), .x8(nXANY), .y9(WSTB));
t391 cell_C15(.x1(NET00121), .x2(NET00122), .y3(NET00121), .y4(NET00119), .x5(IACK), .x6(NET00122), .y9(nV274), .x10(IACK));
t380 cell_D21(.x1(NET00124), .y2(NET00167), .y3(NET00177), .x4(nDIN), .x5(NET00177), .x6(NET00178));
t376 cell_I21(.x1(NET00098), .x3(NET00099), .y4(NET00102), .x6(NET00100), .x8(NET00101), .y9(NET00099));
t376 cell_D16(.x1(NET00101), .x3(NET00031), .y4(NET00089), .x6(NET00089), .x8(NET00114), .y9(NET00090));
t378 cell_J23(.x1(X7), .y2(NET00084), .x3(X6), .x5(nX5));
t416 cell_G17(.c1(NET00145), .q3(NET00034), .d5(C5));
t416 cell_G18(.c1(NET00145), .q4(NET00039), .d5(nC4));
t374 cell_H13(.x1(X2), .x2(NET00008), .x3(X3), .y4(NET00008), .y8(NET00010));
t387 cell_C31(.x1(NET00198), .y2(nCSRRD), .x3(nSYNC), .y4(NET00198), .x5(NET00206), .x6(nCSR));
t381 cell_I27(.x1(X9), .y2(nX6_9), .x3(X8), .x4(X6), .x6(X7));
t390 cell_M27(.x1(NET00022), .y4(Y7IN), .x5(NET00023), .x6(NET00021), .y9(NET00022), .x10(Y7IN));
t416 cell_G20(.c1(NET00145), .q4(NET00100), .d5(nC2));
t377 cell_D27(.x1(NET00041), .y2(NET00172), .x3(NET00101), .y4(NET00173), .x5(nV274), .x6(NET00172), .x8(NET00173), .y9(NET00223));
t406 cell_L27(.c1(X1), .r2(LOCK), .q3(NET00042), .r5(Y7IN), .s10(Y6IN));
t416 cell_G22(.c1(NET00145), .q4(NET00106), .d5(nC0));

endmodule
//______________________________________________________________________________
//
