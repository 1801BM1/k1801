//
// Copyright (c) 2013-2014 by 1801BM1@gmail.com
//______________________________________________________________________________
//
`timescale 1ns / 100ps

module vp_065
(
   inout[15:0] PIN_nAD,       // Address/Data inverted bus
                              //
   input       PIN_nINIT,     //
   input       PIN_nSYNC,     //
   input       PIN_nDIN,      //
   input       PIN_nDOUT,     //
   input       PIN_nBS,       //
   input       PIN_nDCLO,     //
   input       PIN_nIAKI,     //
   output      PIN_nIAKO,     //
   output      PIN_nVIRQ,     //
   output      PIN_nEVNT,     //
   output      PIN_nRPLY,     //
   output      PIN_nSEL,      //
                              //
   output      PIN_nTF,       //
   output      PIN_nRR,       //
   input       PIN_nIP,       //
   input       PIN_nBSYD,     //
                              //
   input       PIN_CLK,       //
   input       PIN_ACL0,      //
   input       PIN_ACL1,      //
   input       PIN_NB0,       //
   input       PIN_NP,        //
   input       PIN_PEV,       //
   input[3:0]  PIN_FR,        //
                              //
   input       GND,           //
   input       VCC            //
);

//______________________________________________________________________________
//
// Autogenerated netlist
//
wire SIM_RESET;

wire nRXCLK;
wire RXIRQ;
wire nTXDATA;
wire TXLD;
wire AD1;
wire n8BIT;
wire nA1;
wire VEC6;
wire nTXTEST;
wire F19200;
wire AD7;
wire TXRDY;
wire PAR;
wire nTXSHC;
wire nTB105;
wire W566;
wire nTCLO;
wire nTXF;
wire AD3;
wire nRXCNT1;
wire R562;
wire nWSTB;
wire TXIER;
wire DIN;
wire nNP;
wire FBAUD;
wire TXTEST;
wire nCLK;
wire TXCNT3;
wire RXLD;
wire TXF;
wire nRXFRAME;
wire nOVFERR;
wire RXLD0;
wire nVECH;
wire VEC2;
wire nRSEL;
wire nA566;
wire R564;
wire W564;
wire PARSET;
wire PARERR;
wire RXFCLR;
wire TXIRQ_ACK;
wire VEC7;
wire nA5;
wire nA3;
wire A566;
wire nRWSEL;
wire nIAKI;
wire nA562;
wire R560;
wire AD0;
wire nFR0;
wire CLK;
wire nSSEL;
wire WSTB;
wire F9600;
wire AD2;
wire n5BIT;
wire TXCNT1;
wire TXCNTL;
wire nTXCNT0B;
wire nTB11;
wire nTXCNT3;
wire NP;
wire nTXCNT0;
wire nTB10;
wire nTXCNT1;
wire nTXCNT2;
wire AD5;
wire AD4;
wire nTB75;
wire nTB12;
wire nTB85;
wire TCLO;
wire TXCNT2;
wire nTB9;
wire TXCNT0;
wire FIX1;
wire n7BIT;
wire nA12;
wire nACL1;
wire TXBRK;
wire RXDIN;
wire AD6;
wire FR0;
wire FR1;
wire nFR1;
wire nTXFRAME;
wire PD8;
wire nTB7;
wire nA2;
wire nBS;
wire nA8;
wire nA10;
wire nFR2;
wire FR2;
wire FR3;
wire nFR3;
wire TXLSB;
wire nA560;
wire nA6;
wire TXSHC;
wire nA4;
wire RXFSET;
wire F57600;
wire nRXEND;
wire nPAR;
wire nA9;
wire A7;
wire nA11;
wire OVFERR;
wire nSYNC;
wire nCLK0;
wire RXIRQ_ACK;
wire TXIRQ;
wire nA564;
wire F150;
wire nF600;
wire F100;
wire F200;
wire RXNEW;
wire F4800;
wire F2400;
wire a8BIT;
wire ITLSB;
wire F1200;
wire DDIN;
wire nRXSTB;
wire TXPCLR;
wire F600;
wire F300;
wire PARCLR;
wire TXSTB;
wire F75;
wire NP0;
wire nRXSTB0;
wire F50;
wire RXBRK;
wire VSEL;
wire TXPSET;
wire TXSTOP;
wire nACL0;
wire nTB6;
wire RXDATA;
wire INIT;
wire RXIER;
wire IRQ_ACK;
wire DOUT;
wire nDIN;
wire RXCLK;
wire VEC3;
wire RXF;
wire RXFRAME;
wire RXSTRT;
wire nRXCNT2;
wire nRXCNT3;
wire RXCNT3;
wire nRXCNT0;
wire nRXSTOP;
wire RXSTB;
wire PD7;
wire nSEL0;
wire TXFRAME;

wire NET00001;
wire NET00003;
wire NET00005;
wire NET00006;
wire NET00007;
wire NET00009;
wire NET00010;
wire NET00035;
wire NET00012;
wire NET00015;
wire NET00017;
wire NET00024;
wire NET00026;
wire NET00028;
wire NET00031;
wire NET00033;
wire NET00034;
wire NET00037;
wire NET00681;
wire NET00038;
wire NET00039;
wire NET00060;
wire NET00040;
wire NET00042;
wire NET00043;
wire NET00046;
wire NET00047;
wire NET00048;
wire NET00022;
wire NET00054;
wire NET00055;
wire NET00056;
wire NET00011;
wire NET00061;
wire NET00062;
wire NET00063;
wire NET00052;
wire NET00064;
wire NET00066;
wire NET00067;
wire NET00459;
wire NET00070;
wire NET00071;
wire NET00072;
wire NET00073;
wire NET00074;
wire NET00075;
wire NET00076;
wire NET00078;
wire NET00079;
wire NET00080;
wire NET00462;
wire NET00084;
wire NET00087;
wire NET00090;
wire NET00091;
wire NET00092;
wire NET00093;
wire NET00095;
wire NET00168;
wire NET00104;
wire NET00105;
wire NET00106;
wire NET00108;
wire NET00111;
wire NET00113;
wire NET00115;
wire NET00116;
wire NET00117;
wire NET00119;
wire NET00122;
wire NET00123;
wire NET00124;
wire NET00126;
wire NET00127;
wire NET00128;
wire NET00136;
wire NET00130;
wire NET00131;
wire NET00133;
wire NET00134;
wire NET00137;
wire NET00415;
wire NET00138;
wire NET00163;
wire NET00143;
wire NET00144;
wire NET00145;
wire NET00146;
wire NET00147;
wire NET00148;
wire NET00149;
wire NET00150;
wire NET00151;
wire NET00153;
wire NET00154;
wire NET00455;
wire NET00156;
wire NET00157;
wire NET00158;
wire NET00172;
wire NET00160;
wire NET00161;
wire NET00162;
wire NET00237;
wire NET00233;
wire NET00165;
wire NET00290;
wire NET00294;
wire NET00351;
wire NET00170;
wire NET00238;
wire NET00234;
wire NET00291;
wire NET00175;
wire NET00176;
wire NET00177;
wire NET00178;
wire NET00179;
wire NET00180;
wire NET00295;
wire NET00182;
wire NET00346;
wire NET00246;
wire NET00487;
wire NET00186;
wire NET00188;
wire NET00194;
wire NET00195;
wire NET00314;
wire NET00359;
wire NET00198;
wire NET00199;
wire NET00200;
wire NET00203;
wire NET00206;
wire NET00207;
wire NET00208;
wire NET00209;
wire NET00210;
wire NET00212;
wire NET00213;
wire NET00303;
wire NET00215;
wire NET00216;
wire NET00219;
wire NET00217;
wire NET00347;
wire NET00463;
wire NET00220;
wire NET00228;
wire NET00222;
wire NET00223;
wire NET00230;
wire NET00225;
wire NET00226;
wire NET00227;
wire NET00480;
wire NET00229;
wire NET00247;
wire NET00231;
wire NET00457;
wire NET00464;
wire NET00488;
wire NET00461;
wire NET00489;
wire NET00456;
wire NET00458;
wire NET00241;
wire NET00245;
wire NET00243;
wire NET00557;
wire NET00517;
wire NET00515;
wire NET00749;
wire NET00250;
wire NET00255;
wire NET00256;
wire NET00257;
wire NET00258;
wire NET00261;
wire NET00264;
wire NET00265;
wire NET00266;
wire NET00267;
wire NET00268;
wire NET00269;
wire NET00273;
wire NET00274;
wire NET00275;
wire NET00276;
wire NET00277;
wire NET00483;
wire NET00279;
wire NET00360;
wire NET00281;
wire NET00301;
wire NET00283;
wire NET00284;
wire NET00285;
wire NET00287;
wire NET00299;
wire NET00289;
wire NET00348;
wire NET00352;
wire NET00362;
wire NET00296;
wire NET00298;
wire NET00358;
wire NET00486;
wire NET00345;
wire NET00772;
wire NET00771;
wire NET00305;
wire NET00307;
wire NET00308;
wire NET00309;
wire NET00310;
wire NET00312;
wire NET00313;
wire NET00315;
wire NET00316;
wire NET00317;
wire NET00318;
wire NET00319;
wire NET00320;
wire NET00699;
wire NET00322;
wire NET00323;
wire NET00324;
wire NET00328;
wire NET00329;
wire NET00330;
wire NET00333;
wire NET00334;
wire NET00336;
wire NET00338;
wire NET00339;
wire NET00340;
wire NET00341;
wire NET00342;
wire NET00343;
wire NET00344;
wire NET00173;
wire NET00414;
wire NET00371;
wire NET00372;
wire NET00349;
wire NET00368;
wire NET00370;
wire NET00594;
wire NET00596;
wire NET00597;
wire NET00598;
wire NET00595;
wire NET00470;
wire NET00472;
wire NET00468;
wire NET00465;
wire NET00471;
wire NET00363;
wire NET00364;
wire NET00021;
wire NET00367;
wire NET00755;
wire NET00752;
wire NET00580;
wire NET00581;
wire NET00579;
wire NET00607;
wire NET00374;
wire NET00606;
wire NET00376;
wire NET00377;
wire NET00380;
wire NET00381;
wire NET00382;
wire NET00384;
wire NET00386;
wire NET00387;
wire NET00390;
wire NET00392;
wire NET00394;
wire NET00395;
wire NET00396;
wire NET00399;
wire NET00400;
wire NET00401;
wire NET00403;
wire NET00801;
wire NET00407;
wire NET00408;
wire NET00409;
wire NET00411;
wire NET00412;
wire NET00413;
wire NET00800;
wire NET00416;
wire NET00417;
wire NET00612;
wire NET00420;
wire NET00421;
wire NET00422;
wire NET00423;
wire NET00424;
wire NET00425;
wire NET00428;
wire NET00429;
wire NET00430;
wire NET00431;
wire NET00434;
wire NET00435;
wire NET00437;
wire NET00438;
wire NET00439;
wire NET00440;
wire NET00441;
wire NET00442;
wire NET00443;
wire NET00444;
wire NET00445;
wire NET00446;
wire NET00447;
wire NET00448;
wire NET00449;
wire NET00450;
wire NET00451;
wire NET00452;
wire NET00453;
wire NET00454;
wire NET00805;
wire NET00799;
wire NET00795;
wire NET00794;
wire NET00798;
wire NET00793;
wire NET00785;
wire NET00786;
wire NET00792;
wire NET00784;
wire NET00779;
wire NET00776;
wire NET00773;
wire NET00473;
wire NET00774;
wire NET00476;
wire NET00479;
wire NET00700;
wire NET00481;
wire NET00775;
wire NET00777;
wire NET00778;
wire NET00627;
wire NET00691;
wire NET00632;
wire NET00633;
wire NET00629;
wire NET00492;
wire NET00493;
wire NET00690;
wire NET00495;
wire NET00496;
wire NET00497;
wire NET00498;
wire NET00501;
wire NET00503;
wire NET00505;
wire NET00506;
wire NET00507;
wire NET00508;
wire NET00509;
wire NET00510;
wire NET00512;
wire NET00513;
wire NET00639;
wire NET00640;
wire NET00643;
wire NET00647;
wire NET00650;
wire NET00648;
wire NET00521;
wire NET00522;
wire NET00645;
wire NET00524;
wire NET00525;
wire NET00637;
wire NET00527;
wire NET00528;
wire NET00529;
wire NET00530;
wire NET00533;
wire NET00534;
wire NET00535;
wire NET00536;
wire NET00538;
wire NET00539;
wire NET00540;
wire NET00541;
wire NET00542;
wire NET00543;
wire NET00544;
wire NET00545;
wire NET00546;
wire NET00547;
wire NET00549;
wire NET00551;
wire NET00552;
wire NET00553;
wire NET00554;
wire NET00555;
wire NET00668;
wire NET00559;
wire NET00560;
wire NET00561;
wire NET00563;
wire NET00564;
wire NET00565;
wire NET00706;
wire NET00567;
wire NET00568;
wire NET00569;
wire NET00686;
wire NET00571;
wire NET00572;
wire NET00573;
wire NET00709;
wire NET00575;
wire NET00576;
wire NET00577;
wire NET00707;
wire NET00705;
wire NET00685;
wire NET00683;
wire NET00582;
wire NET00583;
wire NET00584;
wire NET00585;
wire NET00586;
wire NET00587;
wire NET00682;
wire NET00667;
wire NET00676;
wire NET00671;
wire NET00662;
wire NET00593;
wire NET00669;
wire NET00710;
wire NET00684;
wire NET00708;
wire NET00670;
wire NET00761;
wire NET00758;
wire NET00762;
wire NET00602;
wire NET00760;
wire NET00759;
wire NET00768;
wire NET00769;
wire NET00711;
wire NET00680;
wire NET00610;
wire NET00611;
wire NET00613;
wire NET00614;
wire NET00615;
wire NET00616;
wire NET00617;
wire NET00620;
wire NET00780;
wire NET00621;
wire NET00622;
wire NET00623;
wire NET00624;
wire NET00625;
wire NET00824;
wire NET00765;
wire NET00766;
wire NET00630;
wire NET00764;
wire NET00783;
wire NET00634;
wire NET00807;
wire NET00636;
wire NET00806;
wire NET00825;
wire NET00804;
wire NET00802;
wire NET00641;
wire NET00797;
wire NET00796;
wire NET00782;
wire NET00763;
wire NET00787;
wire NET00651;
wire NET00652;
wire NET00653;
wire NET00654;
wire NET00655;
wire NET00656;
wire NET00657;
wire NET00658;
wire NET00659;
wire NET00788;
wire NET00790;
wire NET00789;
wire NET00729;
wire NET00664;
wire NET00745;
wire NET00838;
wire NET00835;
wire NET00837;
wire NET00821;
wire NET00822;
wire NET00747;
wire NET00744;
wire NET00695;
wire NET00696;
wire NET00694;
wire NET00818;
wire NET00817;
wire NET00678;
wire NET00679;
wire NET00697;
wire NET00698;
wire NET00701;
wire NET00704;
wire NET00808;
wire NET00703;
wire NET00712;
wire NET00713;
wire NET00714;
wire NET00715;
wire NET00719;
wire NET00720;
wire NET00721;
wire NET00724;
wire NET00725;
wire NET00726;
wire NET00810;
wire NET00730;
wire NET00840;
wire NET00731;
wire NET00733;
wire NET00735;
wire NET00736;
wire NET00738;
wire NET00739;
wire NET00740;
wire NET00741;
wire NET00742;
wire NET00743;
wire NET00746;
wire NET00748;
wire NET00751;
wire NET00809;
wire NET00263;
wire NET00812;
wire NET00813;
wire NET00815;
wire NET00816;
wire NET00828;
wire NET00823;
wire NET00829;
wire NET00830;
wire NET00831;
wire NET00832;
wire NET00833;
wire NET00836;

//______________________________________________________________________________
//
// Duplicated cell for power reinforcement
//
// t429 cell_E23(.y3(nRXCLK), .x5(nRXSTB));
// t428 cell_K1(.x2(NET00134), .y3(nCLK));
//

//______________________________________________________________________________
//
// Autogenerated cell instantiations
//
tINPUT cell_PIN9( .y2(AD0),      .x1(PIN_nAD[0]));
tINPUT cell_PIN10(.y2(AD1),      .x1(PIN_nAD[1]));
tINPUT cell_PIN11(.y2(AD2),      .x1(PIN_nAD[2]));
tINPUT cell_PIN12(.y2(AD3),      .x1(PIN_nAD[3]));
tINPUT cell_PIN13(.y2(AD4),      .x1(PIN_nAD[4]));
tINPUT cell_PIN14(.y2(AD5),      .x1(PIN_nAD[5]));
tINPUT cell_PIN15(.y2(AD6),      .x1(PIN_nAD[6]));
tINPUT cell_PIN16(.y2(AD7),      .x1(PIN_nAD[7]));
tINPUT cell_PIN17(.y2(NET00594), .x1(PIN_nAD[8]));
tINPUT cell_PIN18(.y2(NET00597), .x1(PIN_nAD[9]));
tINPUT cell_PIN19(.y2(NET00035), .x1(PIN_nAD[10]));
tINPUT cell_PIN20(.y2(NET00367), .x1(PIN_nAD[11]));
tINPUT cell_PIN22(.y2(NET00370), .x1(PIN_nAD[12]));

tOUTPUT_OE cell_PINOU9( .x1(NET00048), .x2(NET00106), .y1(PIN_nAD[0]));
tOUTPUT_OE cell_PINOU10(.x1(NET00226), .x2(NET00106), .y1(PIN_nAD[1]));
tOUTPUT_OE cell_PINOU11(.x1(NET00342), .x2(NET00106), .y1(PIN_nAD[2]));
tOUTPUT_OE cell_PINOU12(.x1(NET00090), .x2(NET00333), .y1(PIN_nAD[3]));
tOUTPUT_OE cell_PINOU13(.x1(NET00128), .x2(NET00333), .y1(PIN_nAD[4]));
tOUTPUT_OE cell_PINOU14(.x1(NET00126), .x2(NET00333), .y1(PIN_nAD[5]));
tOUTPUT_OE cell_PINOU15(.x1(NET00123), .x2(NET00333), .y1(PIN_nAD[6]));
tOUTPUT_OE cell_PINOU16(.x1(NET00340), .x2(NET00333), .y1(PIN_nAD[7]));
tOUTPUT_OE cell_PINOU22(.x1(NET00527), .x2(NET00106), .y1(PIN_nAD[12]));
tOUTPUT_OE cell_PINOU25(.x1(NET00423), .x2(NET00106), .y1(PIN_nAD[15]));
//
// Simulating unused data bus pins (read-as-zero, write-ignored)
//
tOUTPUT_OE cell_PINOU_8(.x1(1'b1), .x2(NET00106 | NET00333), .y1(PIN_nAD[8]));
tOUTPUT_OE cell_PINOU_9(.x1(1'b1), .x2(NET00106 | NET00333), .y1(PIN_nAD[9]));
tOUTPUT_OE cell_PINOU_10(.x1(1'b1), .x2(NET00106 | NET00333), .y1(PIN_nAD[10]));
tOUTPUT_OE cell_PINOU_11(.x1(1'b1), .x2(NET00106 | NET00333), .y1(PIN_nAD[11]));
tOUTPUT_OE cell_PINOU_13(.x1(1'b1), .x2(NET00106 | NET00333), .y1(PIN_nAD[13]));
tOUTPUT_OE cell_PINOU_14(.x1(1'b1), .x2(NET00106 | NET00333), .y1(PIN_nAD[14]));

tINPUT cell_PIN7( .y2(NET00012), .x1(PIN_NB0));
tINPUT cell_PIN23(.y2(nACL0),    .x1(PIN_ACL0));
tINPUT cell_PIN24(.y2(nACL1),    .x1(PIN_ACL1));
tINPUT cell_PIN30(.y2(nNP),      .x1(PIN_NP));
tINPUT cell_PIN32(.y2(NET00144), .x1(PIN_PEV));
tINPUT cell_PIN3( .y2(nFR0),     .x1(PIN_FR[0]));
tINPUT cell_PIN4( .y2(nFR1),     .x1(PIN_FR[1]));
tINPUT cell_PIN5( .y2(nFR2),     .x1(PIN_FR[2]));
tINPUT cell_PIN6( .y2(nFR3),     .x1(PIN_FR[3]));

tINPUT cell_PIN1( .y2(NET00771), .x1(PIN_CLK));
tINPUT cell_PIN40(.y2(NET00031), .x1(PIN_nDCLO));
tINPUT cell_PIN34(.y2(NET00131), .x1(PIN_nINIT));
tINPUT cell_PIN26(.y2(NET00371), .x1(PIN_nBS));
tINPUT cell_PIN37(.y2(DOUT),     .x1(PIN_nDOUT));
tINPUT cell_PIN38(.y2(NET00147), .x1(PIN_nDIN));
tINPUT cell_PIN41(.y2(NET00414), .x1(PIN_nSYNC));
tINPUT cell_PIN33(.y2(NET00143), .x1(PIN_nIAKI));
tOUTPUT cell_PIN36(.x1(NET00137), .y1(PIN_nIAKO));
tOUTPUT cell_PIN2( .x1(NET00655), .y1(PIN_nEVNT));
tOUTPUT_OC cell_PIN39(.x1(NET00156), .y1(PIN_nRPLY));
tOUTPUT_OC cell_PIN8( .x1(NET00766), .y1(PIN_nSEL));
tOUTPUT_OC cell_PIN35(.x1(NET00136), .y1(PIN_nVIRQ));

tINPUT cell_PIN29(.y2(NET00040), .x1(PIN_nBSYD));
tINPUT cell_PIN28(.y2(NET00454), .x1(PIN_nIP));
tOUTPUT cell_PIN27(.x1(NET00441),.y1(PIN_nTF));
tOUTPUT cell_PIN31(.x1(RXF),     .y1(PIN_nRR));


//______________________________________________________________________________
//
// Refining the initial state for simulation - we should define the flip-flop states
//
assign SIM_RESET = ~PIN_nDCLO;

// t416 cell_O0(.c1(nCLK), .q4(NET00180), .d5(NET00161));
t416 cell_O0(.c1(nCLK), .q4(NET00180), .d5(NET00161 | SIM_RESET));

// t416 cell_O3(.c1(nCLK), .q4(NET00170), .d5(NET00173));
t416 cell_O3(.c1(nCLK), .q4(NET00170), .d5(NET00173 | SIM_RESET));

// t416 cell_O5(.c1(nCLK), .q4(NET00160), .d5(NET00165));
t416 cell_O5(.c1(nCLK), .q4(NET00160), .d5(NET00165 | SIM_RESET));

// t416 cell_O7(.c1(NET00158), .q4(NET00153), .d5(NET00157));
t416 cell_O7(.c1(NET00158 | SIM_RESET), .q4(NET00153), .d5(NET00157 | SIM_RESET));

// t416 cell_O10(.c1(NET00158), .q4(NET00150), .d5(NET00151));
t416 cell_O10(.c1(NET00158 | SIM_RESET), .q4(NET00150), .d5(NET00151 | SIM_RESET));

// t416 cell_N0(.c1(F19200), .q3(NET00800), .q4(NET00801), .d5(NET00799));
t416 cell_N0(.c1(F19200 | SIM_RESET), .q3(NET00800), .q4(NET00801), .d5(NET00799 & ~SIM_RESET));

// t416 cell_N2(.c1(F9600), .q3(NET00794), .q4(NET00795), .d5(NET00793));
t416 cell_N2(.c1(F9600 | SIM_RESET), .q3(NET00794), .q4(NET00795), .d5(NET00793 & ~SIM_RESET));

// t416 cell_N4(.c1(F4800), .q3(NET00785), .q4(NET00786), .d5(NET00784));
t416 cell_N4(.c1(F4800 | SIM_RESET), .q3(NET00785), .q4(NET00786), .d5(NET00784 & ~SIM_RESET));

// t416 cell_N6(.c1(F2400), .q3(NET00777), .q4(NET00778), .d5(NET00776));
t416 cell_N6(.c1(F2400 | SIM_RESET), .q3(NET00777), .q4(NET00778), .d5(NET00776 & ~SIM_RESET));

// t416 cell_N8(.c1(F1200), .q3(NET00773), .q4(NET00774), .d5(nF600));
t416 cell_N8(.c1(F1200 | SIM_RESET), .q3(NET00773), .q4(NET00774), .d5(nF600 & ~SIM_RESET));

// t416 cell_N10(.c1(F600), .q4(NET00690), .d5(NET00632));
t416 cell_N10(.c1(F600 | SIM_RESET), .q4(NET00690), .d5(NET00632 & ~SIM_RESET));

// t416 cell_N11(.c1(nF600), .q3(NET00691), .d5(NET00690));
t416 cell_N11(.c1(nF600 | SIM_RESET), .q3(NET00691), .d5(NET00690 | SIM_RESET));

// t416 cell_L1(.c1(NET00445), .q3(NET00442), .q4(NET00446), .d5(NET00447));
t416 cell_L1(.c1(NET00445 | SIM_RESET), .q3(NET00442), .q4(NET00446), .d5(NET00447 & ~SIM_RESET));

// t416 cell_L3(.c1(NET00450), .q3(NET00448), .q4(NET00451), .d5(NET00452));
t416 cell_L3(.c1(NET00450 | SIM_RESET), .q3(NET00448), .q4(NET00451), .d5(NET00452 & ~SIM_RESET));

// t416 cell_L5(.c1(F150), .q3(NET00430), .q4(NET00434), .d5(NET00435));
t416 cell_L5(.c1(F150 | SIM_RESET), .q3(NET00430), .q4(NET00434), .d5(NET00435 & ~SIM_RESET));

// t416 cell_L7(.c1(F300), .q3(NET00437), .q4(NET00439), .d5(NET00440));
t416 cell_L7(.c1(F300 | SIM_RESET), .q3(NET00437), .q4(NET00439), .d5(NET00440 & ~SIM_RESET));

// t416 cell_L9(.c1(F600), .q3(NET00424), .q4(NET00428), .d5(NET00429));
t416 cell_L9(.c1(F600 | SIM_RESET), .q3(NET00424), .q4(NET00428), .d5(NET00429 & ~SIM_RESET));

// t416 cell_M1(.c1(NET00444), .q3(NET00652), .q4(NET00653), .d5(NET00651));
t416 cell_M1(.c1(NET00444 | SIM_RESET), .q3(NET00652), .q4(NET00653), .d5(NET00651 & ~SIM_RESET));

// t416 cell_M3(.c1(F50), .q3(NET00657), .q4(NET00658), .d5(NET00656));
t416 cell_M3(.c1(F50 | SIM_RESET), .q3(NET00657), .q4(NET00658), .d5(NET00656 & ~SIM_RESET));

// t405 cell_M4(.c1(NET00643), .x2(F100), .q3(F50), .q4(NET00637), .r5(NET00639), .y7(NET00643), .s10(NET00640));
t405 cell_M4(.c1(NET00643 | SIM_RESET ), .x2(F100), .q3(F50), .q4(NET00637), .r5(NET00639), .y7(NET00643), .s10(NET00640));

// t416 cell_M5(.c1(F100), .q3(NET00639), .q4(NET00640), .d5(NET00637));
t416 cell_M5(.c1(F100 | SIM_RESET), .q3(NET00639), .q4(NET00640), .d5(NET00637 & ~SIM_RESET));

// t405 cell_M6(.c1(NET00650), .x2(F200), .q3(F100), .q4(NET00645), .r5(NET00647), .y7(NET00650), .s10(NET00648));
t405 cell_M6(.c1(NET00650 | SIM_RESET), .x2(F200), .q3(F100), .q4(NET00645), .r5(NET00647), .y7(NET00650), .s10(NET00648));

// t416 cell_M7(.c1(F200), .q3(NET00647), .q4(NET00648), .d5(NET00645));
t416 cell_M7(.c1(F200 | SIM_RESET), .q3(NET00647), .q4(NET00648), .d5(NET00645 & ~SIM_RESET));

// t416 cell_M8(.c1(nF600), .q3(NET00632), .q4(NET00633), .d5(NET00629));
t416 cell_M8(.c1(nF600 | SIM_RESET), .q3(NET00632), .q4(NET00633), .d5(NET00629 & ~SIM_RESET));

// t416 cell_M9(.c1(F600), .q4(NET00629), .d5(NET00627));
t416 cell_M9(.c1(F600 | SIM_RESET), .q4(NET00629), .d5(NET00627 & ~SIM_RESET));

// t406 cell_J37(.c1(NET00093), .r2(ITLSB), .q4(TXLSB), .r5(NET00465), .s10(NET00468));
t406 cell_J37(.c1(NET00093 | SIM_RESET), .r2(ITLSB), .q4(TXLSB), .r5(NET00465 | SIM_RESET), .s10(NET00468 & ~SIM_RESET));

// t416 cell_I35(.c1(NET00092), .q4(NET00488), .d5(NET00464));
// t416 cell_H33(.c1(NET00092), .q4(NET00489), .d5(NET00458));
// t416 cell_J27(.c1(NET00092), .q4(NET00186), .d5(NET00179));
// t416 cell_I27(.c1(NET00092), .q4(NET00182), .d5(NET00241));
// t416 cell_I32(.c1(NET00092), .q4(NET00243), .d5(NET00483));
// t416 cell_H30(.c1(NET00092), .q3(NET00517), .d5(NET00360));
// t416 cell_H27(.c1(NET00092), .q4(NET00301), .d5(NET00299));
// t416 cell_G27(.c1(NET00092), .q3(NET00352), .d5(NET00348));
// t406 cell_J36(.c1(NET00471), .r2(ITLSB), .q3(NET00468), .q4(NET00465), .r5(NET00470), .s10(NET00472));
//
t416 cell_I35(.c1(NET00092 | SIM_RESET), .q4(NET00488), .d5(NET00464 | SIM_RESET));
t416 cell_H33(.c1(NET00092 | SIM_RESET), .q4(NET00489), .d5(NET00458 | SIM_RESET));
t416 cell_J27(.c1(NET00092 | SIM_RESET), .q4(NET00186), .d5(NET00179 & ~SIM_RESET));
t416 cell_I27(.c1(NET00092 | SIM_RESET), .q4(NET00182), .d5(NET00241 & ~SIM_RESET));
t416 cell_I32(.c1(NET00092 | SIM_RESET), .q4(NET00243), .d5(NET00483 & ~SIM_RESET));
t416 cell_H30(.c1(NET00092 | SIM_RESET), .q3(NET00517), .d5(NET00360 & ~SIM_RESET));
t416 cell_H27(.c1(NET00092 | SIM_RESET), .q4(NET00301), .d5(NET00299 & ~SIM_RESET));
t416 cell_G27(.c1(NET00092 | SIM_RESET), .q3(NET00352), .d5(NET00348 & ~SIM_RESET));
t406 cell_J36(.c1(NET00471 | SIM_RESET), .r2(ITLSB), .q3(NET00468), .q4(NET00465), .r5(NET00470), .s10(NET00472));

// t405 cell_M30(.c1(NET00070), .x2(NET00070), .q3(TXFRAME), .q4(NET00024), .r5(NET00318), .y7(NET00320), .s10(NET00319));
// t416 cell_M31(.c1(NET00320), .q3(NET00318), .q4(NET00319), .d5(NET00316));
// t416 cell_M25(.c1(FBAUD), .q3(NET00033), .q4(NET00037), .d5(NET00038));
// t405 cell_M26(.c1(NET00034), .x2(FBAUD), .q4(TXRDY), .r5(NET00033), .y7(NET00034), .s10(NET00037));
//
t405 cell_M30(.c1(NET00070 | SIM_RESET), .x2(NET00070), .q3(TXFRAME), .q4(NET00024), .r5(NET00318 | SIM_RESET), .y7(NET00320), .s10(NET00319 & ~SIM_RESET));
t416 cell_M31(.c1(NET00320 | SIM_RESET), .q3(NET00318), .q4(NET00319), .d5(NET00316 & ~SIM_RESET));
t416 cell_M25(.c1(FBAUD | SIM_RESET), .q3(NET00033), .q4(NET00037), .d5(NET00038 & ~SIM_RESET));
t405 cell_M26(.c1(NET00034 | SIM_RESET), .x2(FBAUD), .q4(TXRDY), .r5(NET00033 | SIM_RESET), .y7(NET00034), .s10(NET00037 & ~SIM_RESET));

//______________________________________________________________________________
//
t381 cell_D5(.x1(nSSEL), .y2(NET00407), .x3(DIN), .x4(nWSTB), .x6(nA560));
t370 cell_N26(.y2(NET00829), .x5(nTXCNT0B));
t384 cell_D37(.x1(RXDATA), .y3(RXSTRT), .x5(nRXFRAME));
t429 cell_K19(.y3(nCLK0), .x5(NET00751));
t372 cell_A5(.x1(AD7), .y2(NET00596), .y3(NET00595), .y4(NET00598), .x5(NET00594), .x6(NET00597));
t372 cell_A1(.x1(AD4), .y2(NET00580), .y3(NET00579), .y4(NET00581), .x5(AD5), .x6(AD6));
t428 cell_K4(.x2(NET00145), .y3(W566));
t405 cell_A18(.c1(NET00381), .x2(nRXCLK), .q3(NET00334), .r5(NET00380), .y7(NET00381), .s10(NET00382));
t429 cell_K30(.y3(NET00146), .x5(TXLD));
t406 cell_B6(.c1(nSYNC), .r2(INIT), .q4(nA1), .r5(NET00755), .s10(AD1));
t406 cell_B5(.c1(nSYNC), .r2(INIT), .q4(nA2), .r5(NET00021), .s10(AD2));
t428 cell_E20(.x2(NET00395), .y3(RXNEW));
t428 cell_K21(.x2(NET00080), .y3(NET00113));
t428 cell_K31(.x2(NET00364), .y3(NET00411));
t416 cell_L16(.c1(nCLK), .q3(NET00079), .q4(NET00736), .d5(NET00735));
t384 cell_L14(.x1(DIN), .y3(NET00735), .x5(R562));
t405 cell_A20(.c1(NET00569), .x2(nRXCLK), .q3(NET00528), .r5(NET00567), .y7(NET00569), .s10(NET00568));
t416 cell_A19(.c1(nRXCLK), .q3(NET00380), .q4(NET00382), .d5(NET00279));
t373 cell_B23(.x1(n5BIT), .x3(NET00533), .y4(NET00529));
t384 cell_B22(.x1(OVFERR), .y3(NET00527), .x5(R560));
t388 cell_B9(.x1(NET00322), .y2(NET00760), .x3(nA9), .y4(NET00759), .y5(NET00762), .x6(NET00322), .x7(NET00762), .x10(nA9));
t377 cell_B8(.x1(NET00759), .y2(NET00274), .x3(NET00760), .y4(NET00761), .x5(NET00758), .x6(NET00330), .x8(NET00761), .y9(NET00758));
t406 cell_O28(.c1(NET00810), .r2(nTXFRAME), .q3(TXCNTL), .q4(NET00808), .r5(TXCNT0), .s10(nTXCNT0));
t375 cell_N27(.x1(nTXCNT0B), .y2(NET00206), .y3(NET00810), .x4(NET00263), .x5(NET00263), .x6(TXSHC), .y9(NET00263));
t416 cell_C15(.c1(RXLD0), .q4(NET00283), .d5(NET00281));
t406 cell_O22(.c1(NET00411), .r2(nTXFRAME), .q3(NET00822), .q4(NET00821), .r5(NET00815), .s10(NET00823));
t405 cell_A22(.c1(NET00565), .x2(nRXCLK), .q3(NET00277), .r5(NET00563), .y7(NET00565), .s10(NET00564));
t416 cell_A21(.c1(nRXCLK), .q3(NET00567), .q4(NET00568), .d5(NET00277));
t380 cell_B11(.x1(nA10), .y2(NET00275), .y3(NET00324), .x4(nA11), .x5(NET00324), .x6(nA12));
t405 cell_O23(.c1(NET00812), .x2(NET00411), .q3(NET00815), .q4(NET00823), .r5(NET00821), .y7(NET00812), .s10(NET00822));
t379 cell_C13(.x1(nACL0), .y2(NET00266), .x3(nACL1), .y4(NET00267), .x5(nBS), .x6(nACL0), .x8(nACL1));
t428 cell_E37(.x2(NET00634), .y3(nRXFRAME));
t405 cell_A24(.c1(NET00577), .x2(nRXCLK), .q3(NET00534), .r5(NET00575), .y7(NET00577), .s10(NET00576));
t416 cell_A23(.c1(nRXCLK), .q3(NET00563), .q4(NET00564), .d5(NET00281));
t428 cell_E39(.x2(NET00664), .y3(RXDATA));
t370 cell_D28(.y2(NET00473), .x5(AD6));
t380 cell_N29(.x1(TXCNT1), .y2(nTB105), .y3(NET00828), .x4(NET00829), .x5(NET00828), .x6(nTXCNT3));
t406 cell_O34(.c1(NET00194), .r2(nTXFRAME), .q3(NET00195), .q4(NET00198), .r5(TXCNT3), .s10(nTXCNT3));
t406 cell_A29(.c1(NET00582), .r2(NET00546), .q3(NET00583), .q4(NET00585), .r5(NET00507), .s10(NET00584));
t416 cell_B21(.c1(NET00339), .q4(NET00336), .d5(NET00376));
t384 cell_L24(.x1(FBAUD), .y3(NET00070), .x5(NET00026));
t416 cell_A25(.c1(nRXCLK), .q3(NET00575), .q4(NET00576), .d5(RXDIN));
t416 cell_B17(.c1(RXLD0), .q4(NET00087), .d5(NET00289));
t416 cell_B16(.c1(RXLD0), .q4(NET00127), .d5(NET00334));
t373 cell_L25(.x1(W566), .x3(nCLK0), .y4(NET00063));
t380 cell_N31(.x1(nTXCNT0B), .y2(nTB11), .y3(NET00258), .x4(nTXCNT1), .x5(NET00258), .x6(nTXCNT3));
t387 cell_M29(.x1(NET00024), .y2(NET00026), .x3(TXFRAME), .y4(TXLD), .x5(TXRDY), .x6(TXRDY));
t405 cell_O27(.c1(NET00818), .x2(NET00816), .q3(TXSHC), .q4(NET00074), .r5(NET00817), .y7(NET00818), .s10(NET00052));
t406 cell_O26(.c1(NET00816), .r2(nTXFRAME), .q3(NET00052), .q4(NET00817), .r5(TXSHC), .s10(NET00074));
t416 cell_B19(.c1(nRXCLK), .q3(NET00343), .q4(NET00344), .d5(NET00334));
t405 cell_B18(.c1(NET00349), .x2(nRXCLK), .q3(NET00289), .r5(NET00343), .y7(NET00349), .s10(NET00344));
t374 cell_B27(.x1(nNP), .x2(RXDATA), .x3(NET00541), .y4(NET00539), .y8(NET00541));
t372 cell_B4(.x1(AD1), .y2(NET00021), .y3(NET00755), .y4(NET00752), .x5(AD2), .x6(AD3));
t393 cell_B26(.x1(NET00538), .x3(NET00539), .y4(NET00540), .x5(nNP), .x6(NET00540), .y9(RXDIN));
t416 cell_L26(.c1(NET00061), .q3(NET00067), .d5(NET00066));
t416 cell_L27(.c1(NET00063), .q4(NET00066), .d5(NET00062));
t393 cell_B20(.x1(NET00528), .x3(NET00529), .y4(NET00530), .x5(n5BIT), .x6(NET00530), .y9(NET00279));
t384 cell_L30(.x1(TXFRAME), .y3(NET00363), .x5(nTCLO));
t406 cell_A2(.c1(nSYNC), .r2(INIT), .q4(nA5), .r5(NET00580), .s10(AD5));
t416 cell_C17(.c1(RXLD0), .q4(NET00124), .d5(NET00279));
t416 cell_C16(.c1(RXLD0), .q4(NET00054), .d5(NET00277));
t373 cell_L31(.x1(FBAUD), .x3(NET00363), .y4(NET00364));
t417 cell_D10(.x1(R562), .y4(NET00047), .x5(NET00222), .x6(NET00055), .x10(TXBRK));
t404 cell_A34(.c1(nRXCNT0), .q3(NET00741), .q4(nRXCNT1), .r5(NET00748), .s10(NET00749));
t406 cell_A4(.c1(nSYNC), .r2(INIT), .q3(A7), .r5(NET00595), .s10(AD7));
t384 cell_D11(.x1(R562), .y3(NET00226), .x5(NET00225));
t416 cell_C19(.c1(nRXCLK), .q3(NET00284), .q4(NET00287), .d5(NET00289));
t375 cell_B25(.x1(NET00533), .y2(NET00535), .y3(a8BIT), .x4(a8BIT), .x5(n8BIT), .x6(RXDIN), .y9(NET00533));
t393 cell_B24(.x1(NET00534), .x3(NET00535), .y4(NET00536), .x5(a8BIT), .x6(NET00536), .y9(NET00281));
t406 cell_B29(.c1(NET00507), .r2(NET00546), .q3(NET00544), .q4(NET00542), .r5(NET00508), .s10(NET00545));
t406 cell_A7(.c1(nSYNC), .r2(INIT), .q4(nA9), .r5(NET00598), .s10(NET00597));
t405 cell_C18(.c1(NET00285), .x2(nRXCLK), .q3(NET00217), .r5(NET00284), .y7(NET00285), .s10(NET00287));
t405 cell_C21(.c1(NET00493), .x2(nRXCLK), .q3(NET00223), .r5(NET00492), .y7(NET00493), .s10(NET00495));
t416 cell_C20(.c1(nRXCLK), .q3(NET00492), .q4(NET00495), .d5(NET00217));
t405 cell_C23(.c1(NET00497), .x2(nRXCLK), .q3(NET00220), .r5(NET00496), .y7(NET00497), .s10(NET00498));
t405 cell_B28(.c1(NET00543), .x2(NET00507), .q3(NET00508), .q4(NET00545), .r5(NET00542), .y7(NET00543), .s10(NET00544));
t405 cell_L28(.c1(NET00061), .x2(NET00063), .q3(NET00062), .r5(NET00060), .y7(NET00061), .s10(NET00064));
t416 cell_L29(.c1(NET00063), .q3(NET00060), .q4(NET00064), .d5(TXLD));
t406 cell_A10(.c1(nSYNC), .r2(INIT), .q4(nA11), .r5(NET00607), .s10(NET00367));
t371 cell_A9(.x1(NET00035), .y3(NET00606), .y4(NET00607), .x6(NET00367));
t381 cell_L33(.x1(n7BIT), .y2(NET00313), .x3(nTB9), .x4(NP), .x6(FIX1));
t381 cell_L34(.x1(n7BIT), .y2(NET00312), .x3(nTB9), .x4(nNP), .x6(GND));
t416 cell_C22(.c1(nRXCLK), .q3(NET00496), .q4(NET00498), .d5(NET00223));
t384 cell_C37(.x1(RXSTRT), .y3(NET00704), .x5(nRXSTOP));
t371 cell_A12(.x1(NET00370), .y3(NET00368), .y4(NET00372), .x6(NET00371));
t406 cell_A11(.c1(nSYNC), .r2(INIT), .q4(nA12), .r5(NET00368), .s10(NET00370));
t406 cell_B31(.c1(NET00508), .r2(NET00546), .q3(NET00712), .q4(NET00714), .r5(NET00510), .s10(NET00713));
t405 cell_B30(.c1(NET00715), .x2(NET00508), .q3(NET00510), .q4(NET00713), .r5(NET00714), .y7(NET00715), .s10(NET00712));
t390 cell_M23(.x1(nTXF), .y4(NET00039), .x5(NET00040), .x6(nTCLO), .y9(NET00038), .x10(NET00039));
t406 cell_N24(.c1(NET00813), .r2(nTXFRAME), .q3(NET00830), .q4(NET00832), .r5(NET00816), .s10(NET00831));
t383 cell_B2(.x1(nA4), .y2(NET00273), .x3(nA5), .x4(nA6), .x5(A7), .x6(nA8));
t406 cell_B1(.c1(nSYNC), .r2(INIT), .q4(nA4), .r5(NET00579), .s10(AD4));
t381 cell_L35(.x1(n7BIT), .y2(NET00310), .x3(nTB10), .x4(nNP), .x6(FIX1));
t406 cell_A13(.c1(nSYNC), .r2(INIT), .q4(nBS), .r5(NET00372), .s10(NET00371));
t381 cell_L36(.x1(n8BIT), .y2(NET00308), .x3(nTB12), .x4(NP), .x6(GND));
t381 cell_O38(.x1(nTXCNT2), .y2(NET00188), .x3(TXCNTL), .x4(nTXCNT1), .x6(nTXCNT0));
t380 cell_O37(.x1(nTXCNT2), .y2(nTB7), .y3(NET00203), .x4(nTXCNT1), .x5(NET00203), .x6(nTXCNT0));
t376 cell_B33(.x1(nRXCNT0), .x3(nRXCNT3), .y4(NET00719), .x6(nRXCNT1), .x8(nRXCNT3), .y9(NET00720));
t417 cell_D12(.x1(R562), .y4(NET00227), .x5(NET00219), .x6(NET00055), .x10(TXTEST));
t417 cell_B32(.x1(nNP), .y4(NET00698), .x5(NET00720), .x6(NP0), .x10(NET00719));
t391 cell_C7(.x1(nA2), .x2(nA2), .y3(NET00111), .y4(nA560), .x5(nA1), .x6(NET00111), .y9(nA564), .x10(nA1));
t373 cell_G33(.x1(TXSTB), .x3(NET00525), .y4(NET00559));
t387 cell_B12(.x1(nACL0), .y2(NET00322), .x3(nA3), .y4(NET00323), .x5(nACL1), .x6(nACL1));
t388 cell_B10(.x1(NET00329), .y2(NET00329), .x3(NET00323), .y4(NET00330), .y5(NET00328), .x6(nA3), .x7(NET00328), .x10(nACL1));
t383 cell_O25(.x1(NET00074), .y2(TXSTB), .x3(NET00813), .x4(NET00816), .x5(NET00812), .x6(NET00815));
t373 cell_C1(.x1(NET00106), .x3(nVECH), .y4(NET00108));
t406 cell_D26(.c1(NET00407), .r2(INIT), .q3(RXIER), .r5(NET00473), .s10(AD6));
t388 cell_C9(.x1(nA1), .y2(NET00119), .x3(nA2), .y4(A566), .y5(nA562), .x6(NET00119), .x7(nA1), .x10(nA2));
t381 cell_L38(.x1(n8BIT), .y2(NET00307), .x3(nTB11), .x4(nNP), .x6(GND));
t404 cell_A32(.c1(nRXCNT1), .q3(NET00739), .q4(nRXCNT2), .r5(NET00738), .s10(NET00740));
t370 cell_O39(.y2(nTB75), .x5(NET00188));
t376 cell_C24(.x1(PARSET), .x3(NET00503), .y4(NET00392), .x6(NET00505), .x8(PARCLR), .y9(NET00390));
t416 cell_H34(.c1(nCLK0), .q3(NET00525), .d5(NET00524));
t406 cell_A8(.c1(nSYNC), .r2(INIT), .q4(nA10), .r5(NET00606), .s10(NET00035));
t406 cell_A6(.c1(nSYNC), .r2(INIT), .q4(nA8), .r5(NET00596), .s10(NET00594));
t406 cell_A3(.c1(nSYNC), .r2(INIT), .q4(nA6), .r5(NET00581), .s10(AD6));
t386 cell_D7(.x1(NET00408), .y2(NET00408), .y3(nSEL0), .y4(NET00409), .x5(NET00269), .x6(nSYNC), .x7(VCC));
t370 cell_D23(.y2(nRXSTB), .x5(RXSTB));
t394 cell_C12(.x1(NET00265), .y2(NET00265), .x3(NET00266), .y4(NET00268), .x5(NET00264), .x6(NET00268), .y9(NET00269), .x10(NET00267));
t373 cell_D31(.x1(FBAUD), .x3(NET00546), .y4(NET00636));
t385 cell_D29(.x1(nNP), .x2(NET00401), .y3(NET00401), .x5(NET00400), .y8(NET00403));
t406 cell_B3(.c1(nSYNC), .r2(INIT), .q4(nA3), .r5(NET00752), .s10(AD3));
t381 cell_G36(.x1(nTXFRAME), .y2(TXPSET), .x3(TXLSB), .x4(NET00552), .x6(NET00551));
t405 cell_O29(.c1(NET00809), .x2(NET00810), .q3(TXCNT0), .q4(nTXCNT0), .r5(NET00808), .y7(NET00809), .s10(TXCNTL));
t376 cell_C33(.x1(n7BIT), .x3(NET00697), .y4(NET00699), .x6(n8BIT), .x8(NET00698), .y9(NET00700));
t428 cell_E36(.x2(NET00630), .y3(DDIN));
t373 cell_F15(.x1(NET00084), .x3(nRXEND), .y4(RXLD));
t370 cell_H2(.y2(nDIN), .x5(DIN));
t376 cell_I19(.x1(NET00064), .x3(NET00067), .y4(ITLSB), .x6(NET00031), .x8(ITLSB), .y9(NET00001));
t416 cell_A15(.c1(nCLK), .q4(NET00376), .d5(NET00374));
t370 cell_F36(.y2(NET00554), .x5(NET00144));
t376 cell_H39(.x1(n8BIT), .x3(nTB10), .y4(NET00512), .x6(n7BIT), .x8(nTB105), .y9(NET00513));
t405 cell_O31(.c1(NET00210), .x2(NET00206), .q3(TXCNT1), .q4(NET00208), .r5(NET00209), .y7(NET00210), .s10(NET00207));
t416 cell_H26(.c1(NET00093), .q4(NET00298), .d5(NET00296));
t376 cell_H25(.x1(NET00298), .x3(NET00115), .y4(NET00303), .x6(NET00295), .x8(NET00303), .y9(NET00299));
t375 cell_D36(.x1(NET00113), .y2(NET00679), .y3(NET00678), .x4(INIT), .x5(INIT), .x6(NET00679), .y9(NET00630));
t373 cell_H21(.x1(NET00294), .x3(NET00117), .y4(NET00295));
t429 cell_K2(.y3(F57600), .x5(NET00133));
t384 cell_D22(.x1(nRXFRAME), .y3(NET00476), .x5(RXDATA));
t417 cell_G5(.x1(R562), .y4(NET00128), .x5(NET00127), .x6(VSEL), .x10(VCC));
t385 cell_F7(.x1(NET00764), .x2(NET00765), .y3(NET00765), .x5(NET00409), .y8(NET00766));
t391 cell_F2(.x1(VSEL), .x2(NET00768), .y3(NET00342), .y4(NET00769), .x5(VEC2), .x6(NET00769), .y9(NET00768), .x10(NET00227));
t417 cell_H38(.x1(NET00512), .y4(NET00840), .x5(nNP), .x6(NET00513), .x10(nNP));
t416 cell_G23(.c1(W566), .q3(NET00351), .d5(AD7));
t416 cell_G21(.c1(W566), .q3(NET00294), .d5(AD6));
t428 cell_K0(.x2(NET00138), .y3(CLK));
t374 cell_G28(.x1(NET00352), .x2(a8BIT), .x3(NET00362), .y4(NET00296), .y8(NET00362));
t383 cell_C29(.x1(NET00507), .y2(RXSTB), .x3(NET00508), .x4(NET00510), .x5(NET00506), .x6(NET00509));
t416 cell_J3(.c1(VCC), .q3(NET00154), .q4(NET00158), .d5(F57600));
t373 cell_I23(.x1(NET00237), .x3(NET00117), .y4(NET00238));
t416 cell_I21(.c1(W566), .q3(NET00237), .d5(AD3));
t416 cell_A16(.c1(NET00339), .q4(NET00374), .d5(NET00377));
t416 cell_A27(.c1(nRXCLK), .q3(NET00571), .q4(NET00572), .d5(RXDATA));
t417 cell_F10(.x1(R562), .y4(NET00090), .x5(NET00087), .x6(VSEL), .x10(VEC3));
t406 cell_G15(.c1(W564), .r2(INIT), .q3(TXBRK), .r5(NET00042), .s10(AD0));
t416 cell_H37(.c1(nCLK0), .q4(NET00521), .d5(TXSTOP));
t404 cell_A28(.c1(NET00509), .q3(NET00507), .q4(NET00584), .r5(NET00585), .s10(NET00583));
t416 cell_G30(.c1(NET00093), .q4(NET00358), .d5(NET00301));
t416 cell_J22(.c1(W566), .q3(NET00168), .d5(AD1));
t373 cell_F21(.x1(NET00394), .x3(NET00384), .y4(NET00395));
t417 cell_H6(.x1(R562), .y4(NET00422), .x5(NET00283), .x6(NET00055), .x10(TXF));
t416 cell_A39(.c1(NET00009), .q3(nOVFERR), .q4(OVFERR), .d5(NET00726));
t373 cell_G24(.x1(NET00351), .x3(NET00117), .y4(NET00346));
t385 cell_H15(.x1(NET00012), .x2(GND), .y3(n7BIT), .x5(n5BIT), .y8(n5BIT));
t416 cell_G26(.c1(NET00093), .q4(NET00345), .d5(GND));
t373 cell_H29(.x1(NET00290), .x3(NET00117), .y4(NET00291));
t429 cell_E1(.y3(NET00333), .x5(NET00108));
t384 cell_A38(.x1(NET00582), .y3(NET00509), .x5(VCC));
t406 cell_H17(.c1(W564), .r2(INIT), .q3(TXIER), .r5(NET00017), .s10(AD6));
t416 cell_H23(.c1(W566), .q3(NET00290), .d5(AD5));
t402 cell_F33(.r1(NET00559), .q3(NET00602), .s6(nTXFRAME));
t416 cell_F22(.c1(NET00011), .q4(NET00394), .d5(NET00396));
t370 cell_H35(.y2(NET00522), .x5(nCLK0));
t428 cell_E3(.x2(NET00105), .y3(VSEL));
t380 cell_A14(.x1(NET00104), .y2(NET00341), .y3(nVECH), .x4(nACL0), .x5(nACL0), .x6(nACL1));
t428 cell_E5(.x2(NET00412), .y3(R562));
t406 cell_I17(.c1(nCLK), .r2(nRWSEL), .q3(NET00782), .q4(NET00156), .r5(GND), .s10(NET00797));
t378 cell_F38(.x1(NET00611), .y2(NET00441), .x3(TCLO), .x5(NET00610));
t406 cell_A35(.c1(NET00746), .r2(nRXFRAME), .q3(NET00749), .q4(NET00748), .r5(NET00741), .s10(nRXCNT1));
t428 cell_E6(.x2(NET00116), .y3(R560));
t405 cell_L17(.c1(NET00731), .x2(nCLK), .q3(NET00733), .r5(NET00079), .y7(NET00731), .s10(NET00736));
t428 cell_E29(.x2(NET00453), .y3(RXFRAME));
t381 cell_L39(.x1(n8BIT), .y2(NET00309), .x3(nTB9), .x4(nNP), .x6(FIX1));
t374 cell_F39(.x1(nTXDATA), .x2(NET00040), .x3(TXBRK), .y4(NET00611), .y8(NET00610));
t376 cell_G25(.x1(NET00345), .x3(NET00115), .y4(NET00347), .x6(NET00346), .x8(NET00347), .y9(NET00348));
t379 cell_F27(.x1(nPAR), .y2(PAR), .x3(NET00390), .y4(nPAR), .x5(RXNEW), .x6(NET00392), .x8(PAR));
t371 cell_B35(.x1(nRXCNT0), .y3(NET00721), .y4(NET00479), .x6(NET00721));
t399 cell_H18(.r1(W566), .x2(NET00001), .q3(TXF), .q4(nTXF), .s6(NET00003), .y7(NET00003));
t428 cell_E7(.x2(NET00409), .y3(nSSEL));
t417 cell_B34(.x1(nNP), .y4(NET00697), .x5(NET00719), .x6(NP0), .x10(RXCNT3));
t377 cell_J0(.x1(NET00772), .y2(NET00772), .x3(CLK), .y4(NET00134), .x5(NET00771), .x6(nCLK), .x8(NET00771), .y9(NET00138));
t373 cell_J8(.x1(RXIRQ), .x3(TXIRQ), .y4(NET00136));
t405 cell_F25(.c1(NET00011), .x2(nCLK0), .q3(NET00386), .r5(NET00384), .y7(NET00011), .s10(NET00387));
t428 cell_E15(.x2(RXLD), .y3(RXLD0));
t406 cell_O30(.c1(NET00206), .r2(nTXFRAME), .q3(NET00207), .q4(NET00209), .r5(TXCNT1), .s10(NET00208));
t405 cell_M2(.c1(NET00659), .x2(F50), .q3(NET00450), .q4(NET00656), .r5(NET00657), .y7(NET00659), .s10(NET00658));
t391 cell_H3(.x1(R560), .x2(NET00420), .y3(NET00340), .y4(NET00423), .x5(PARERR), .x6(NET00422), .y9(NET00420), .x10(NET00421));
t405 cell_O33(.c1(NET00216), .x2(NET00212), .q3(TXCNT2), .q4(nTXCNT2), .r5(NET00215), .y7(NET00216), .s10(NET00213));
t405 cell_L0(.c1(NET00443), .x2(NET00445), .q3(NET00444), .q4(NET00447), .r5(NET00442), .y7(NET00443), .s10(NET00446));
t406 cell_O32(.c1(NET00212), .r2(nTXFRAME), .q3(NET00213), .q4(NET00215), .r5(TXCNT2), .s10(nTXCNT2));
t429 cell_E22(.y3(nRXCLK), .x5(nRXSTB));
t405 cell_L4(.c1(NET00431), .x2(F150), .q3(F75), .q4(NET00435), .r5(NET00430), .y7(NET00431), .s10(NET00434));
t405 cell_O35(.c1(NET00199), .x2(NET00194), .q3(TXCNT3), .q4(nTXCNT3), .r5(NET00198), .y7(NET00199), .s10(NET00195));
t405 cell_N1(.c1(NET00805), .x2(F19200), .q3(F9600), .q4(NET00799), .r5(NET00800), .y7(NET00805), .s10(NET00801));
t416 cell_O1(.c1(CLK), .q3(NET00176), .d5(NET00180));
t372 cell_G17(.x1(AD0), .y2(NET00043), .y3(NET00042), .y4(NET00017), .x5(AD2), .x6(AD6));
t372 cell_L22(.x1(NET00072), .y2(NET00072), .y3(NET00073), .y4(NET00071), .x5(NET00071), .x6(NET00074));
t377 cell_O2(.x1(NET00162), .y2(NET00133), .x3(NET00176), .y4(NET00173), .x5(NET00175), .x6(NET00162), .x8(NET00160), .y9(NET00175));
t405 cell_N3(.c1(NET00798), .x2(F9600), .q3(F4800), .q4(NET00793), .r5(NET00794), .y7(NET00798), .s10(NET00795));
t405 cell_M0(.c1(NET00654), .x2(NET00444), .q3(NET00655), .q4(NET00651), .r5(NET00652), .y7(NET00654), .s10(NET00653));
t405 cell_L2(.c1(NET00449), .x2(NET00450), .q3(NET00445), .q4(NET00452), .r5(NET00448), .y7(NET00449), .s10(NET00451));
t406 cell_F20(.c1(RXNEW), .r2(INIT), .q3(RXBRK), .r5(NET00229), .s10(NET00231));
t389 cell_M32(.x1(NET00315), .x2(NET00317), .y3(NET00316), .x4(TCLO), .y5(NET00315), .x6(PD8), .x10(PD7));
t373 cell_D39(.x1(nRXEND), .x3(OVFERR), .y4(NET00006));
t428 cell_K35(.x2(NET00363), .y3(nTXFRAME));
t417 cell_H5(.x1(VSEL), .y4(NET00421), .x5(VEC7), .x6(R560), .x10(RXF));
t417 cell_G6(.x1(R562), .y4(NET00126), .x5(NET00124), .x6(VSEL), .x10(VCC));
t387 cell_B14(.x1(nACL1), .y2(VEC7), .x3(NET00341), .y4(VEC3), .x5(nACL0), .x6(nACL1));
t417 cell_G10(.x1(NET00054), .y4(NET00056), .x5(R562), .x6(NET00055), .x10(TXIER));
t385 cell_G7(.x1(VEC6), .x2(NET00122), .y3(NET00122), .x5(NET00056), .y8(NET00123));
t385 cell_H14(.x1(n5BIT), .x2(NET00012), .y3(n8BIT), .x5(NET00015), .y8(NET00015));
t389 cell_F32(.x1(TXLSB), .x2(NET00593), .y3(TXPCLR), .x4(NET00551), .y5(NET00551), .x6(TXSTB), .x10(NET00602));
t416 cell_H32(.c1(NET00093), .q4(NET00486), .d5(NET00515));
t374 cell_G32(.x1(NET00517), .x2(n5BIT), .x3(NET00557), .y4(NET00515), .y8(NET00557));
t376 cell_G29(.x1(NET00358), .x3(NET00115), .y4(NET00359), .x6(NET00291), .x8(NET00359), .y9(NET00360));
t373 cell_J23(.x1(NET00163), .x3(NET00117), .y4(NET00172));
t416 cell_J21(.c1(W566), .q3(NET00163), .d5(AD2));
t428 cell_E4(.x2(R564), .y3(NET00055));
t428 cell_E2(.x2(NET00134), .y3(nCLK));
t406 cell_G18(.c1(W564), .r2(INIT), .q3(TXTEST), .q4(nTXTEST), .r5(NET00043), .s10(AD2));
t418 cell_F28(.x1(NET00399), .x2(NET00144), .y3(NET00399), .y4(NET00400), .x5(nPAR), .x6(NET00144), .x10(PAR));
t379 cell_F37(.x1(NET00593), .y2(NET00552), .x3(NET00586), .y4(NET00593), .x5(nTXFRAME), .x6(NET00587), .x8(NET00552));
t406 cell_N22(.c1(NET00815), .r2(nTXFRAME), .q3(NET00835), .q4(NET00837), .r5(NET00813), .s10(NET00836));
t393 cell_G14(.x1(R560), .x3(NET00046), .y4(NET00048), .x5(RXBRK), .x6(NET00047), .y9(NET00046));
t416 cell_J9(.c1(nDIN), .q3(NET00612), .q4(NET00614), .d5(TXIRQ));
t376 cell_I30(.x1(NET00486), .x3(NET00115), .y4(NET00487), .x6(NET00234), .x8(NET00487), .y9(NET00483));
t373 cell_I29(.x1(NET00233), .x3(NET00117), .y4(NET00234));
t428 cell_K14(.x2(NET00763), .y3(WSTB));
t405 cell_N5(.c1(NET00792), .x2(F4800), .q3(F2400), .q4(NET00784), .r5(NET00785), .y7(NET00792), .s10(NET00786));
t428 cell_K12(.x2(NET00711), .y3(FBAUD));
t416 cell_I33(.c1(NET00093), .q4(NET00456), .d5(NET00186));
t428 cell_K15(.x2(NET00147), .y3(DIN));
t416 cell_I28(.c1(W566), .q3(NET00233), .d5(AD4));
t416 cell_O8(.c1(NET00154), .q3(NET00149), .d5(NET00153));
t405 cell_N9(.c1(NET00775), .x2(F1200), .q3(F600), .q4(nF600), .r5(NET00773), .y7(NET00775), .s10(NET00774));
t384 cell_J28(.x1(nTXSHC), .y3(NET00091), .x5(NET00146));
t374 cell_J12(.x1(NET00782), .x2(DOUT), .x3(NET00783), .y4(NET00763), .y8(NET00783));
t429 cell_K5(.y3(nIAKI), .x5(NET00143));
t406 cell_I9(.c1(DIN), .r2(INIT), .q3(NET00613), .q4(NET00615), .r5(NET00612), .s10(NET00614));
t376 cell_O9(.x1(NET00148), .x3(NET00149), .y4(NET00151), .x6(NET00148), .x8(NET00150), .y9(F19200));
t405 cell_L6(.c1(NET00438), .x2(F300), .q3(F150), .q4(NET00440), .r5(NET00437), .y7(NET00438), .s10(NET00439));
t374 cell_J7(.x1(TXIRQ_ACK), .x2(NET00764), .x3(RXIRQ_ACK), .y4(NET00764), .y8(IRQ_ACK));
t376 cell_M10(.x1(NET00633), .x3(NET00691), .y4(NET00627), .x6(NET00633), .x8(NET00629), .y9(F200));
t388 cell_I12(.x1(NET00824), .y2(NET00788), .x3(NET00789), .y4(TXIRQ), .y5(NET00824), .x6(TXF), .x7(NET00824), .x10(TXIER));
t406 cell_I11(.c1(NET00824), .r2(TXIRQ_ACK), .q3(NET00787), .q4(NET00790), .r5(GND), .s10(VCC));
t383 cell_L11(.x1(F150), .y2(NET00706), .x3(nFR0), .x4(nFR1), .x5(FR2), .x6(FR3));
t376 cell_J25(.x1(NET00177), .x3(NET00115), .y4(NET00178), .x6(NET00172), .x8(NET00178), .y9(NET00179));
t376 cell_I25(.x1(NET00245), .x3(NET00115), .y4(NET00246), .x6(NET00238), .x8(NET00246), .y9(NET00241));
t405 cell_N7(.c1(NET00779), .x2(F2400), .q3(F1200), .q4(NET00776), .r5(NET00777), .y7(NET00779), .s10(NET00778));
t416 cell_I26(.c1(NET00093), .q4(NET00245), .d5(NET00243));
t416 cell_O6(.c1(CLK), .q3(NET00161), .q4(NET00162), .d5(NET00160));
t405 cell_I15(.c1(NET00825), .x2(nCLK), .q3(NET00802), .r5(NET00806), .y7(NET00825), .s10(NET00807));
t377 cell_I7(.x1(NET00625), .y2(NET00137), .x3(NET00613), .y4(NET00624), .x5(NET00624), .x6(NET00625), .x8(NET00615), .y9(TXIRQ_ACK));
t406 cell_J11(.c1(NET00788), .r2(INIT), .q3(NET00789), .r5(NET00787), .s10(NET00790));
t405 cell_L8(.c1(NET00425), .x2(F600), .q3(F300), .q4(NET00429), .r5(NET00424), .y7(NET00425), .s10(NET00428));
t416 cell_I3(.c1(nDIN), .q3(NET00620), .q4(NET00621), .d5(RXIRQ));
t416 cell_O4(.c1(CLK), .q4(NET00165), .d5(NET00170));
t428 cell_K6(.x2(NET00413), .y3(W564));
t416 cell_J26(.c1(NET00093), .q4(NET00177), .d5(NET00182));
t416 cell_O11(.c1(NET00154), .q3(NET00157), .q4(NET00148), .d5(NET00150));
t406 cell_I5(.c1(DIN), .r2(INIT), .q3(NET00622), .q4(NET00623), .r5(NET00620), .s10(NET00621));
t416 cell_I16(.c1(NET00825), .q4(NET00796), .d5(NET00804));
t370 cell_I37(.y2(NET00471), .x5(NET00093));
t403 cell_J13(.x1(NET00269), .x2(nRSEL), .x3(IRQ_ACK), .y4(nRSEL), .x5(DIN), .x6(NET00269), .y7(NET00780), .x8(NET00780), .y9(nRWSEL), .x10(DOUT));
t416 cell_J16(.c1(nCLK), .q4(NET00804), .d5(NET00802));
t405 cell_N23(.c1(NET00838), .x2(NET00815), .q3(NET00813), .q4(NET00836), .r5(NET00837), .y7(NET00838), .s10(NET00835));
t416 cell_I34(.c1(NET00093), .q4(NET00461), .d5(NET00489));
t416 cell_I36(.c1(NET00093), .q3(NET00472), .q4(NET00470), .d5(NET00488));
t405 cell_A36(.c1(NET00745), .x2(RXCLK), .q3(NET00746), .q4(nRXCNT0), .r5(NET00744), .y7(NET00745), .s10(NET00747));
t416 cell_J15(.c1(nCLK), .q3(NET00806), .q4(NET00807), .d5(nRWSEL));
t373 cell_J17(.x1(nRWSEL), .x3(NET00796), .y4(NET00797));
t383 cell_O16(.x1(F2400), .y2(NET00667), .x3(FR0), .x4(FR1), .x5(FR2), .x6(nFR3));
t383 cell_N16(.x1(F200), .y2(NET00686), .x3(FR0), .x4(FR1), .x5(nFR2), .x6(FR3));
t406 cell_A37(.c1(RXCLK), .r2(nRXFRAME), .q3(NET00747), .q4(NET00744), .r5(NET00746), .s10(nRXCNT0));
t381 cell_M34(.x1(NET00310), .y2(PD7), .x3(NET00312), .x4(NET00314), .x6(NET00313));
t428 cell_K20(.x2(nRSEL), .y3(NET00106));
t406 cell_C31(.c1(NET00510), .r2(NET00546), .q3(NET00696), .q4(NET00694), .r5(NET00641), .s10(NET00506));
t428 cell_K23(.x2(TXLD), .y3(NET00115));
t429 cell_K24(.y3(NET00117), .x5(TXLD));
t373 cell_J34(.x1(NET00459), .x3(NET00117), .y4(NET00462));
t376 cell_J35(.x1(NET00461), .x3(NET00115), .y4(NET00463), .x6(NET00462), .x8(NET00463), .y9(NET00464));
t371 cell_N12(.x1(nFR2), .y3(FR2), .y4(FR3), .x6(nFR3));
t371 cell_O12(.x1(nFR0), .y3(FR0), .y4(FR1), .x6(nFR1));
t383 cell_N13(.x1(F1200), .y2(NET00685), .x3(nFR0), .x4(nFR1), .x5(nFR2), .x6(FR3));
t373 cell_J30(.x1(NET00168), .x3(NET00117), .y4(NET00455));
t416 cell_J32(.c1(W566), .q3(NET00459), .d5(AD0));
t383 cell_M12(.x1(F100), .y2(NET00709), .x3(FR0), .x4(nFR1), .x5(FR2), .x6(FR3));
t387 cell_M16(.x1(NET00708), .y2(NET00710), .x3(NET00710), .y4(NET00711), .x5(NET00684), .x6(NET00670));
t383 cell_O13(.x1(F19200), .y2(NET00671), .x3(nFR0), .x4(nFR1), .x5(FR2), .x6(nFR3));
t383 cell_N14(.x1(F600), .y2(NET00683), .x3(FR0), .x4(nFR1), .x5(nFR2), .x6(FR3));
t405 cell_C30(.c1(NET00695), .x2(NET00510), .q3(NET00641), .q4(NET00506), .r5(NET00694), .y7(NET00695), .s10(NET00696));
t383 cell_O15(.x1(F4800), .y2(NET00676), .x3(nFR0), .x4(FR1), .x5(FR2), .x6(nFR3));
t383 cell_N15(.x1(F300), .y2(NET00682), .x3(nFR0), .x4(FR1), .x5(nFR2), .x6(FR3));
t383 cell_M15(.x1(NET00705), .y2(NET00708), .x3(NET00707), .x4(NET00709), .x5(NET00706), .x6(NET00686));
t376 cell_J33(.x1(NET00456), .x3(NET00115), .y4(NET00457), .x6(NET00455), .x8(NET00457), .y9(NET00458));
t383 cell_M13(.x1(F75), .y2(NET00707), .x3(nFR0), .x4(FR1), .x5(FR2), .x6(FR3));
t383 cell_O14(.x1(F9600), .y2(NET00669), .x3(FR0), .x4(nFR1), .x5(FR2), .x6(nFR3));
t383 cell_M14(.x1(F50), .y2(NET00705), .x3(FR0), .x4(FR1), .x5(FR2), .x6(FR3));
t428 cell_K28(.x2(nTXSHC), .y3(NET00093));
t428 cell_K29(.x2(NET00091), .y3(NET00092));
t381 cell_M38(.x1(n5BIT), .y2(NET00257), .x3(nTB75), .x4(nNP), .x6(GND));
t381 cell_M39(.x1(n5BIT), .y2(NET00255), .x3(nTB85), .x4(NP), .x6(GND));
t379 cell_C34(.x1(NET00701), .y2(nRXSTOP), .x3(NET00699), .y4(NET00701), .x5(NET00700), .x6(n5BIT), .x8(NET00703));
t429 cell_K37(.y3(nSYNC), .x5(NET00414));
t428 cell_K38(.x2(NET00131), .y3(INIT));
t405 cell_M27(.c1(nCLK0), .x2(TXF), .q3(TCLO), .q4(nTCLO), .r5(NET00028), .y7(NET00028), .s10(NET00031));
t380 cell_C25(.x1(nRXSTB0), .y2(nRXSTB0), .y3(PARCLR), .x4(nPAR), .x5(RXSTB), .x6(NET00501));
t370 cell_J19(.y2(NET00751), .x5(nCLK));
t383 cell_N17(.x1(NET00682), .y2(NET00684), .x3(NET00683), .x4(NET00685), .x5(NET00667), .x6(NET00676));
t380 cell_O17(.x1(NET00669), .y2(NET00670), .y3(NET00668), .x4(NET00671), .x5(NET00668), .x6(NET00662));
t378 cell_N32(.x1(NET00263), .y2(NET00212), .x3(nTXCNT0B), .x5(nTXCNT1));
t383 cell_O18(.x1(nFR3), .y2(NET00662), .x3(FR0), .x4(FR1), .x5(nFR2), .x6(F57600));
t381 cell_N33(.x1(nTXCNT2), .y2(NET00194), .x3(nTXCNT0B), .x4(nTXCNT1), .x6(NET00263));
t416 cell_L18(.c1(nCLK), .q4(NET00730), .d5(NET00733));
t416 cell_D16(.c1(RXLD0), .q4(NET00225), .d5(NET00223));
t390 cell_N35(.x1(TXCNT1), .y4(nTB9), .x5(TXCNT3), .x6(TXCNT2), .y9(nTB12), .x10(TXCNT3));
t370 cell_N36(.y2(nTXCNT1), .x5(TXCNT1));
t385 cell_D21(.x1(NET00476), .x2(INIT), .y3(NET00230), .x5(NET00480), .y8(NET00480));
t373 cell_L20(.x1(NET00078), .x3(NET00079), .y4(NET00080));
t406 cell_A33(.c1(NET00741), .r2(nRXFRAME), .q3(NET00740), .q4(NET00738), .r5(NET00739), .s10(nRXCNT2));
t374 cell_B15(.x1(NET00336), .x2(nCLK), .x3(NET00338), .y4(NET00130), .y8(NET00339));
t381 cell_N37(.x1(NET00255), .y2(NET00256), .x3(NET00257), .x4(NET00247), .x6(NET00250));
t406 cell_F18(.c1(RXLD0), .r2(DDIN), .q3(RXF), .r5(RXFCLR), .s10(RXFSET));
t404 cell_D18(.c1(RXNEW), .q3(RXFSET), .q4(RXFCLR), .r5(NET00231), .s10(NET00229));
t402 cell_D19(.r1(NET00228), .q3(NET00229), .q4(NET00231), .s6(NET00230));
t406 cell_C39(.c1(NET00006), .r2(DDIN), .q3(NET00007), .q4(NET00010), .r5(NET00005), .s10(NET00009));
t418 cell_B36(.x1(nNP), .x2(nNP), .y3(NP0), .y4(NET00703), .x5(NET00724), .x6(NP0), .x10(NET00725));
t404 cell_A30(.c1(nRXCNT2), .q3(RXCNT3), .q4(nRXCNT3), .r5(NET00742), .s10(NET00743));
t416 cell_F23(.c1(nCLK0), .q4(NET00396), .d5(NET00386));
t387 cell_I39(.x1(nNP), .y2(nTB6), .x3(n5BIT), .y4(NET00481), .x5(NET00481), .x6(NET00022));
t371 cell_C38(.x1(NET00454), .y3(NET00680), .y4(NET00681), .x6(nTXTEST));
t380 cell_O36(.x1(nTXCNT2), .y2(NET00022), .y3(NET00200), .x4(nTXCNT1), .x5(NET00200), .x6(TXCNT0));
t385 cell_G38(.x1(NET00840), .x2(TXSTOP), .y3(TXSTOP), .x5(nTB6), .y8(NET00560));
t374 cell_C2(.x1(IRQ_ACK), .x2(NET00104), .x3(NET00095), .y4(NET00104), .y8(NET00105));
t418 cell_G39(.x1(TXSTOP), .x2(TXLSB), .y3(NET00561), .y4(nTXDATA), .x5(NET00555), .x6(NET00561), .x10(NET00560));
t370 cell_N28(.y2(nTXCNT0B), .x5(TXCNT0));
t428 cell_E32(.x2(NET00641), .y3(RXCLK));
t380 cell_N30(.x1(TXCNT1), .y2(nTB10), .y3(NET00261), .x4(nTXCNT0B), .x5(NET00261), .x6(nTXCNT3));
t381 cell_L32(.x1(n7BIT), .y2(NET00314), .x3(nTB11), .x4(NP), .x6(GND));
t406 cell_C36(.c1(NET00678), .r2(INIT), .q3(NET00453), .q4(NET00634), .r5(NET00704), .s10(RXCLK));
t405 cell_N25(.c1(NET00833), .x2(NET00813), .q3(NET00816), .q4(NET00831), .r5(NET00832), .y7(NET00833), .s10(NET00830));
t405 cell_A26(.c1(NET00573), .x2(nRXCLK), .q3(NET00538), .r5(NET00571), .y7(NET00573), .s10(NET00572));
t381 cell_L37(.x1(n8BIT), .y2(NET00305), .x3(nTB11), .x4(NP), .x6(FIX1));
t416 cell_F17(.c1(RXFRAME), .q4(NET00084), .d5(RXF));
t428 cell_E34(.x2(NET00636), .y3(NET00582));
t429 cell_E14(.y3(nRXEND), .x5(NET00130));
t373 cell_D20(.x1(nRXSTB0), .x3(NET00479), .y4(NET00228));
t379 cell_C27(.x1(NET00503), .y2(NET00505), .x3(PARCLR), .y4(NET00503), .x5(RXNEW), .x6(PARSET), .x8(NET00505));
t379 cell_G34(.x1(NET00547), .y2(NET00549), .x3(TXPCLR), .y4(NET00547), .x5(nTXFRAME), .x6(TXPSET), .x8(NET00549));
t381 cell_D3(.x1(nSSEL), .y2(NET00412), .x3(nSEL0), .x4(WSTB), .x6(nA562));
t406 cell_B39(.c1(NET00005), .r2(DDIN), .q3(NET00726), .r5(OVFERR), .s10(nOVFERR));
t381 cell_C3(.x1(nSSEL), .y2(NET00095), .x3(nSEL0), .x4(WSTB), .x6(nA566));
t381 cell_D2(.x1(nSSEL), .y2(R564), .x3(nSEL0), .x4(WSTB), .x6(nA564));
t416 cell_H36(.c1(NET00522), .q4(NET00524), .d5(NET00521));
t417 cell_D38(.x1(NET00680), .y4(NET00664), .x5(nTXTEST), .x6(NET00681), .x10(nTXDATA));
t372 cell_L23(.x1(NET00076), .y2(NET00076), .y3(nTXSHC), .y4(NET00075), .x5(NET00075), .x6(NET00073));
t370 cell_M33(.y2(NET00317), .x5(NET00256));
t381 cell_M37(.x1(NET00305), .y2(PD8), .x3(NET00307), .x4(NET00309), .x6(NET00308));
t416 cell_D15(.c1(RXLD0), .q4(NET00219), .d5(NET00217));
t416 cell_D17(.c1(RXLD0), .q4(NET00222), .d5(NET00220));
t416 cell_A17(.c1(nCLK), .q3(NET00338), .q4(NET00377), .d5(nRXFRAME));
t384 cell_N34(.x1(TXCNTL), .y3(nTB85), .x5(TXCNT3));
t416 cell_F26(.c1(nCLK0), .q3(NET00384), .q4(NET00387), .d5(RXFRAME));
t379 cell_B37(.x1(nRXCNT2), .y2(NET00724), .x3(nRXCNT1), .y4(NET00725), .x5(nRXCNT0), .x6(nRXCNT2), .x8(nRXCNT1));
t406 cell_F29(.c1(RXLD0), .r2(DDIN), .q3(PARERR), .r5(NET00401), .s10(NET00403));
t416 cell_L19(.c1(NET00731), .q4(NET00078), .d5(NET00730));
t429 cell_E33(.y3(NET00546), .x5(RXSTRT));
t406 cell_A31(.c1(NET00739), .r2(nRXFRAME), .q3(NET00743), .q4(NET00742), .r5(RXCNT3), .s10(nRXCNT3));
t418 cell_G37(.x1(NET00552), .x2(NET00552), .y3(NET00553), .y4(NET00555), .x5(NET00144), .x6(NET00553), .x10(NET00554));
t417 cell_G9(.x1(VSEL), .y4(VEC6), .x5(VEC7), .x6(R560), .x10(RXIER));
t381 cell_C4(.x1(nSSEL), .y2(NET00116), .x3(nSEL0), .x4(WSTB), .x6(nA560));
t388 cell_H0(.x1(NET00415), .y2(NET00417), .x3(NET00416), .y4(RXIRQ), .y5(NET00415), .x6(RXIER), .x7(NET00415), .x10(RXF));
t406 cell_I0(.c1(NET00415), .r2(RXIRQ_ACK), .q3(NET00616), .q4(NET00617), .r5(GND), .s10(VCC));
t377 cell_J5(.x1(nIAKI), .y2(NET00625), .x3(NET00622), .y4(VEC2), .x5(VEC2), .x6(nIAKI), .x8(NET00623), .y9(RXIRQ_ACK));
t406 cell_I1(.c1(NET00417), .r2(INIT), .q3(NET00416), .r5(NET00616), .s10(NET00617));
t382 cell_C10(.x1(NET00274), .y2(NET00264), .x3(NET00275), .x4(NET00276), .x5(NET00273), .x6(nBS), .y8(NET00276));
t382 cell_D8(.x1(nSSEL), .y2(NET00413), .x3(nWSTB), .x4(DIN), .x5(WSTB), .x6(nA564), .y8(nWSTB));
t382 cell_C26(.x1(RXNEW), .y2(PARSET), .x3(NET00501), .x4(PAR), .x5(RXDATA), .x6(nRXSTB0), .y8(NET00501));
t382 cell_N38(.x1(n5BIT), .y2(NET00250), .x3(nTB7), .x4(nNP), .x5(GND), .x6(FIX1), .y8(FIX1));
t382 cell_D4(.x1(nSSEL), .y2(NET00145), .x3(DIN), .x4(nWSTB), .x5(A566), .x6(nA566), .y8(nA566));
t382 cell_N39(.x1(n5BIT), .y2(NET00247), .x3(nTXCNT3), .x4(NP), .x5(nNP), .x6(FIX1), .y8(NP));
t405 cell_B38(.c1(NET00729), .x2(NET00006), .q3(NET00005), .q4(NET00009), .r5(NET00010), .y7(NET00729), .s10(NET00007));
t376 cell_F35(.x1(NET00549), .x3(TXPCLR), .y4(NET00586), .x6(TXPSET), .x8(NET00547), .y9(NET00587));

endmodule
//______________________________________________________________________________
//
