//
// Copyright (c) 2021 by 1801BM1@gmail.com
//______________________________________________________________________________
//
`timescale 1ns / 100ps

module vp_034
(
   input[1:0]  PIN_RC,        // configuration select
   inout[15:0] PIN_nAD,       // Address/Data inverted bus
   input[15:0] PIN_nD,        // Data/Pattern input
                              //
   input       PIN_nDME,      //
   input       PIN_nCA,       //
   input       PIN_nCB,       //
   input       PIN_nCD,       //
   input       PIN_C,         //
   inout       PIN_nCOM       //
);

//______________________________________________________________________________
//
// Autogenerated netlist
//
wire GND = 1'b0;

wire DMEX0;
wire DME1;
wire VIRQ;
wire D9;
wire D10;
wire D11;
wire D12;
wire D13;
wire D14;
wire D15;
wire R2;
wire R5;
wire R9;
wire R10;
wire R13;
wire R14;
wire R12;
wire R11;
wire COM;
wire PD1;
wire PD2;
wire PD3;
wire PD4;
wire AD4;
wire AD5;
wire PD5;
wire AD6;
wire PD6;
wire AD7;
wire PD7;
wire RC1;
wire MATCH;
wire R0;
wire D5;
wire D7;
wire D8;
wire AD3;
wire R15;
wire R8;
wire R4;
wire D2;
wire D1;
wire R7;
wire D4;
wire D3;
wire R6;
wire R3;
wire R1;
wire CB;
wire nAD13;
wire nCA;
wire nRC1;
wire nCB;
wire nRC0;
wire RC3;
wire nDME3;
wire PD0;
wire nCOM;
wire RIRQ;
wire nRC3;
wire RC0;
wire nCD;
wire D0;
wire CA;
wire D6;

wire NET00000;
wire NET00001;
wire NET00002;
wire NET00003;
wire NET00004;
wire NET00005;
wire NET00148;
wire NET00008;
wire NET00009;
wire NET00249;
wire NET00011;
wire NET00012;
wire NET00013;
wire NET00010;
wire NET00262;
wire NET00022;
wire NET00023;
wire NET00024;
wire NET00025;
wire NET00033;
wire NET00254;
wire NET00035;
wire NET00255;
wire NET00252;
wire NET00042;
wire NET00043;
wire NET00044;
wire NET00045;
wire NET00046;
wire NET00047;
wire NET00048;
wire NET00049;
wire NET00050;
wire NET00051;
wire NET00052;
wire NET00053;
wire NET00054;
wire NET00055;
wire NET00056;
wire NET00057;
wire NET00251;
wire NET00060;
wire NET00061;
wire NET00064;
wire NET00065;
wire NET00253;
wire NET00067;
wire NET00068;
wire NET00071;
wire NET00162;
wire NET00073;
wire NET00074;
wire NET00076;
wire NET00166;
wire NET00079;
wire NET00080;
wire NET00083;
wire NET00088;
wire NET00085;
wire NET00100;
wire NET00093;
wire NET00090;
wire NET00186;
wire NET00185;
wire NET00095;
wire NET00098;
wire NET00218;
wire NET00217;
wire NET00219;
wire NET00108;
wire NET00119;
wire NET00241;
wire NET00121;
wire NET00122;
wire NET00123;
wire NET00126;
wire NET00127;
wire NET00128;
wire NET00129;
wire NET00130;
wire NET00131;
wire NET00132;
wire NET00133;
wire NET00134;
wire NET00135;
wire NET00138;
wire NET00139;
wire NET00140;
wire NET00141;
wire NET00142;
wire NET00143;
wire NET00257;
wire NET00146;
wire NET00007;
wire NET00149;
wire NET00259;
wire NET00152;
wire NET00153;
wire NET00154;
wire NET00155;
wire NET00156;
wire NET00158;
wire NET00159;
wire NET00160;
wire NET00161;
wire NET00211;
wire NET00210;
wire NET00164;
wire NET00165;
wire NET00209;
wire NET00167;
wire NET00168;
wire NET00169;
wire NET00170;
wire NET00171;
wire NET00172;
wire NET00174;
wire NET00175;
wire NET00176;
wire NET00178;
wire NET00179;
wire NET00180;
wire NET00181;
wire NET00182;
wire NET00183;
wire NET00238;
wire NET00256;
wire NET00189;
wire NET00190;
wire NET00191;
wire NET00192;
wire NET00236;
wire NET00194;
wire NET00195;
wire NET00196;
wire NET00223;
wire NET00198;
wire NET00199;
wire NET00200;
wire NET00201;
wire NET00202;
wire NET00203;
wire NET00204;
wire NET00205;
wire NET00206;
wire NET00207;
wire NET00208;
wire NET00234;
wire NET00235;
wire NET00233;
wire NET00242;
wire NET00214;
wire NET00215;
wire NET00216;
wire NET00228;
wire NET00232;
wire NET00226;
wire NET00220;
wire NET00222;
wire NET00229;
wire NET00248;
wire NET00224;
wire NET00247;
wire NET00227;
wire NET00244;
wire NET00243;
wire NET00230;
wire NET00245;
wire NET00237;
wire NET00240;
wire NET00239;
wire NET00250;
wire NET00246;
wire NET00260;
wire NET00261;

//______________________________________________________________________________
//
// Autogenerated cell instantiations
//
tINPUT      cell_PIN2(.y1(RC0),       .x1(PIN_RC[0]));
tINPUT      cell_PIN1(.y1(NET00250),  .x1(PIN_RC[1]));

tINPUT      cell_PIN9(. y2(NET00060), .x1(PIN_nAD[0]));
tINPUT      cell_PIN10(.y2(NET00067), .x1(PIN_nAD[1]));
tINPUT      cell_PIN11(.y2(NET00073), .x1(PIN_nAD[2]));
tINPUT      cell_PIN12(.y2(AD3),      .x1(PIN_nAD[3]));
tINPUT      cell_PIN13(.y2(AD4),      .x1(PIN_nAD[4]));
tINPUT      cell_PIN14(.y2(AD5),      .x1(PIN_nAD[5]));
tINPUT      cell_PIN15(.y2(AD6),      .x1(PIN_nAD[6]));
tINPUT      cell_PIN16(.y2(AD7),      .x1(PIN_nAD[7]));
tINPUT      cell_PIN17(.y2(NET00237), .x1(PIN_nAD[8]));
tINPUT      cell_PIN18(.y2(NET00239), .x1(PIN_nAD[9]));
tINPUT      cell_PIN19(.y2(NET00240), .x1(PIN_nAD[10]));
tINPUT      cell_PIN20(.y2(NET00214), .x1(PIN_nAD[11]));
tINPUT      cell_PIN22(.y2(NET00215), .x1(PIN_nAD[12]));
tINPUT      cell_PIN23(.y2(NET00129), .x1(PIN_nAD[13]));

tOUTPUT_OE  cell_PINOU9( .x1(NET00024), .x2(NET00002), .y1(PIN_nAD[0]));
tOUTPUT_OE  cell_PINOU10(.x1(NET00013), .x2(NET00002), .y1(PIN_nAD[1]));
tOUTPUT_OE  cell_PINOU11(.x1(NET00023), .x2(NET00001), .y1(PIN_nAD[2]));
tOUTPUT_OE  cell_PINOU12(.x1(NET00011), .x2(NET00001), .y1(PIN_nAD[3]));
tOUTPUT_OE  cell_PINOU13(.x1(NET00010), .x2(NET00001), .y1(PIN_nAD[4]));
tOUTPUT_OE  cell_PINOU14(.x1(NET00003), .x2(NET00001), .y1(PIN_nAD[5]));
tOUTPUT_OE  cell_PINOU15(.x1(NET00005), .x2(NET00001), .y1(PIN_nAD[6]));
tOUTPUT_OE  cell_PINOU16(.x1(NET00022), .x2(NET00001), .y1(PIN_nAD[7]));
tOUTPUT_OE  cell_PINOU17(.x1(NET00080), .x2(NET00000), .y1(PIN_nAD[8]));
tOUTPUT_OE  cell_PINOU18(.x1(NET00042), .x2(NET00000), .y1(PIN_nAD[9]));
tOUTPUT_OE  cell_PINOU19(.x1(NET00043), .x2(NET00000), .y1(PIN_nAD[10]));
tOUTPUT_OE  cell_PINOU20(.x1(NET00051), .x2(NET00000), .y1(PIN_nAD[11]));
tOUTPUT_OE  cell_PINOU22(.x1(NET00050), .x2(NET00000), .y1(PIN_nAD[12]));
tOUTPUT_OE  cell_PINOU23(.x1(NET00049), .x2(NET00000), .y1(PIN_nAD[13]));
tOUTPUT_OE  cell_PINOU24(.x1(NET00048), .x2(NET00000), .y1(PIN_nAD[14]));
tOUTPUT_OE  cell_PINOU25(.x1(NET00047), .x2(NET00000), .y1(PIN_nAD[15]));

tINPUT      cell_PIN26(.y2(D0),  .x1(PIN_nD[0]));
tINPUT      cell_PIN27(.y2(D1),  .x1(PIN_nD[1]));
tINPUT      cell_PIN28(.y2(D2),  .x1(PIN_nD[2]));
tINPUT      cell_PIN29(.y2(D3),  .x1(PIN_nD[3]));
tINPUT      cell_PIN30(.y2(D4),  .x1(PIN_nD[4]));
tINPUT      cell_PIN31(.y2(D5),  .x1(PIN_nD[5]));
tINPUT      cell_PIN32(.y2(D6),  .x1(PIN_nD[6]));
tINPUT      cell_PIN33(.y2(D7),  .x1(PIN_nD[7]));
tINPUT      cell_PIN3( .y2(D8),  .x1(PIN_nD[8]));
tINPUT      cell_PIN4( .y2(D9),  .x1(PIN_nD[9]));
tINPUT      cell_PIN5( .y2(D10), .x1(PIN_nD[10]));
tINPUT      cell_PIN6( .y2(D11), .x1(PIN_nD[11]));
tINPUT      cell_PIN7( .y2(D12), .x1(PIN_nD[12]));
tINPUT      cell_PIN8( .y2(D13), .x1(PIN_nD[13]));
tINPUT      cell_PIN35(.y2(D14), .x1(PIN_nD[14]));
tINPUT      cell_PIN36(.y2(D15), .x1(PIN_nD[15]));

tINPUT      cell_PIN34(.y1(NET00174), .x1(PIN_nDME));
tINPUT      cell_PIN41(.y1(NET00153), .x1(PIN_nCA));
tINPUT      cell_PIN38(.y1(NET00176), .x1(PIN_nCB));
tINPUT      cell_PIN37(.y1(NET00175), .x1(PIN_nCD));
tINPUT      cell_PIN39(.y2(NET00155), .x1(PIN_nCOM));
tINPUT      cell_PIN40(.y1(NET00149), .x1(PIN_C));

tOUTPUT_OE  cell_PINOU39(.x1(nDME3), .x2(NET00180), .y1(PIN_nCOM));

//______________________________________________________________________________
//
t420 cell_A0(.x1(R5), .y2(NET00003), .y3(NET00004), .x4(NET00004), .x5(DMEX0), .x6(NET00223), .x7(NET00233), .x10(NET00007));
t420 cell_A2(.x1(R6), .y2(NET00005), .y3(NET00008), .x4(NET00008), .x5(DMEX0), .x6(NET00192), .x7(NET00235), .x10(NET00007));
t420 cell_D0(.x1(R3), .y2(NET00011), .y3(NET00012), .x4(NET00012), .x5(DMEX0), .x6(NET00143), .x7(NET00207), .x10(NET00007));
t420 cell_C0(.x1(R4), .y2(NET00010), .y3(NET00009), .x4(NET00009), .x5(DMEX0), .x6(NET00160), .x7(NET00161), .x10(NET00007));
t419 cell_G0(.x1(R1), .y2(NET00013), .x4(VIRQ), .x5(DMEX0), .x6(NET00170), .x10(NET00007));
t416 cell_M0(.c1(NET00035), .q4(R13), .d5(D13));
t416 cell_N0(.c1(NET00035), .q4(R11), .d5(D11));
t416 cell_O0(.c1(NET00035), .q4(R9), .d5(D9));
t419 cell_I0(.x1(R0), .y2(NET00024), .x4(MATCH), .x5(DMEX0), .x6(NET00229), .x10(NET00007));
t416 cell_M1(.c1(NET00035), .q4(R12), .d5(D12));
t416 cell_N1(.c1(NET00035), .q4(R10), .d5(D10));
t416 cell_O1(.c1(NET00035), .q4(R8), .d5(D8));
t420 cell_F0(.x1(R2), .y2(NET00023), .y3(NET00033), .x4(NET00033), .x5(DMEX0), .x6(NET00196), .x7(NET00242), .x10(NET00007));
t420 cell_A3(.x1(R7), .y2(NET00022), .y3(NET00025), .x4(NET00025), .x5(DMEX0), .x6(NET00122), .x7(NET00234), .x10(NET00007));
t392 cell_A16(.x1(R10), .x3(NET00046), .y4(NET00043), .x5(NET00044));
t392 cell_A24(.x1(R12), .x3(NET00053), .y4(NET00050), .x5(NET00044));
t392 cell_A32(.x1(R14), .x3(NET00055), .y4(NET00048), .x5(NET00044));
t392 cell_A12(.x1(R9), .x3(NET00045), .y4(NET00042), .x5(NET00044));
t392 cell_A20(.x1(R11), .x3(NET00052), .y4(NET00051), .x5(NET00044));
t392 cell_A28(.x1(R13), .x3(NET00054), .y4(NET00049), .x5(NET00044));
t392 cell_A36(.x1(R15), .x3(NET00056), .y4(NET00047), .x5(NET00044));
t406 cell_C29(.c1(NET00057), .r2(DME1), .q4(NET00093), .r5(NET00219), .s10(AD6));
t395 cell_C4(.x1(PD0), .y2(NET00064), .x3(NET00064), .x4(nCOM), .x5(nCOM), .x6(PD0), .y8(NET00065));
t395 cell_C32(.x1(PD7), .y2(NET00098), .x3(NET00098), .x4(nCOM), .x5(nCOM), .x6(PD7), .y8(NET00056));
t395 cell_C8(.x1(PD1), .y2(NET00262), .x3(NET00262), .x4(nCOM), .x5(nCOM), .x6(PD1), .y8(NET00045));
t392 cell_A8(.x1(R8), .x3(NET00065), .y4(NET00080), .x5(NET00044));
t395 cell_C12(.x1(PD2), .y2(NET00071), .x3(NET00071), .x4(nCOM), .x5(nCOM), .x6(PD2), .y8(NET00046));
t395 cell_C16(.x1(PD3), .y2(NET00076), .x3(NET00076), .x4(nCOM), .x5(nCOM), .x6(PD3), .y8(NET00052));
t395 cell_C20(.x1(PD4), .y2(NET00085), .x3(NET00085), .x4(nCOM), .x5(nCOM), .x6(PD4), .y8(NET00053));
t395 cell_C24(.x1(PD5), .y2(NET00090), .x3(NET00090), .x4(nCOM), .x5(nCOM), .x6(PD5), .y8(NET00054));
t395 cell_C28(.x1(PD6), .y2(NET00095), .x3(NET00095), .x4(nCOM), .x5(nCOM), .x6(PD6), .y8(NET00055));
t406 cell_C33(.c1(NET00057), .r2(DME1), .q4(NET00100), .r5(NET00241), .s10(AD7));
t406 cell_C5(.c1(NET00057), .r2(DME1), .q4(NET00061), .r5(NET00162), .s10(NET00060));
t406 cell_C9(.c1(NET00057), .r2(DME1), .q4(NET00068), .r5(NET00166), .s10(NET00067));
t406 cell_C13(.c1(NET00057), .r2(DME1), .q4(NET00074), .r5(NET00186), .s10(NET00073));
t406 cell_C17(.c1(NET00057), .r2(DME1), .q4(NET00079), .r5(NET00185), .s10(AD3));
t406 cell_C21(.c1(NET00057), .r2(DME1), .q4(NET00083), .r5(NET00218), .s10(AD4));
t406 cell_C25(.c1(NET00057), .r2(DME1), .q4(NET00088), .r5(NET00217), .s10(AD5));
t374 cell_D17(.x1(NET00079), .x2(AD3), .x3(nCD), .y4(PD3), .y8(NET00185));
t429 cell_E32(.y3(nCD), .x5(NET00199));
t395 cell_G6(.x1(D4), .y2(NET00168), .x3(NET00168), .x4(AD7), .x5(AD7), .x6(D4), .y8(NET00169));
t395 cell_I6(.x1(D15), .y2(NET00238), .x3(NET00238), .x4(NET00215), .x5(NET00215), .x6(D15), .y8(NET00211));
t381 cell_I28(.x1(RC3), .y2(NET00189), .x3(NET00044), .x4(CB), .x6(CA));
t372 cell_L18(.x1(NET00244), .y2(NET00244), .y3(NET00245), .y4(NET00243), .x5(NET00243), .x6(NET00246));
t374 cell_D25(.x1(NET00088), .x2(AD5), .x3(nCD), .y4(PD5), .y8(NET00217));
t395 cell_G10(.x1(D2), .y2(NET00140), .x3(NET00140), .x4(AD5), .x5(AD5), .x6(D2), .y8(NET00131));
t372 cell_J5(.x1(NET00255), .y2(NET00255), .y3(NET00002), .y4(NET00254), .x5(NET00254), .x6(NET00253));
t371 cell_J35(.x1(NET00216), .y3(NET00208), .y4(NET00216), .x6(DMEX0));
t374 cell_D29(.x1(NET00093), .x2(AD6), .x3(nCD), .y4(PD6), .y8(NET00219));
t374 cell_D33(.x1(NET00100), .x2(AD7), .x3(nCD), .y4(PD7), .y8(NET00241));
t395 cell_G14(.x1(D0), .y2(NET00138), .x3(NET00138), .x4(AD3), .x5(AD3), .x6(D0), .y8(NET00132));
t416 cell_H7(.c1(nCA), .q4(MATCH), .d5(NET00126));
t429 cell_K10(.y3(nRC1), .x5(NET00250));
t374 cell_D21(.x1(NET00083), .x2(AD4), .x3(nCD), .y4(PD4), .y8(NET00218));
t417 cell_G19(.x1(D3), .y4(NET00141), .x5(CA), .x6(D11), .x10(CB));
t417 cell_H19(.x1(D7), .y4(NET00119), .x5(CA), .x6(D15), .x10(CB));
t372 cell_O32(.x1(NET00183), .y2(NET00183), .y3(NET00181), .y4(NET00182), .x5(NET00182), .x6(nDME3));
t428 cell_K34(.x2(NET00208), .y3(NET00044));
t429 cell_K33(.y3(NET00108), .x5(NET00146));
t372 cell_L17(.x1(NET00248), .y2(NET00248), .y3(NET00249), .y4(NET00247), .x5(NET00247), .x6(NET00245));
t372 cell_F21(.x1(NET00206), .y2(NET00206), .y3(NET00204), .y4(NET00205), .x5(NET00205), .x6(NET00159));
t429 cell_K23(.y3(NET00165), .x5(nDME3));
t417 cell_G25(.x1(D2), .y4(NET00194), .x5(CA), .x6(D10), .x10(CB));
t390 cell_M17(.x1(D8), .y4(NET00242), .x5(NET00165), .x6(D9), .y9(NET00207), .x10(NET00165));
t428 cell_K35(.x2(NET00198), .y3(DMEX0));
t376 cell_L20(.x1(NET00158), .x3(DMEX0), .y4(NET00159), .x6(nRC0), .x8(RC1), .y9(NET00158));
t428 cell_K26(.x2(NET00152), .y3(CA));
t389 cell_L29(.x1(nRC0), .x2(NET00149), .y3(NET00148), .x4(RC1), .y5(NET00146), .x6(NET00149), .x10(nRC0));
t378 cell_L31(.x1(RC1), .y2(NET00200), .x3(NET00176), .x5(nRC0));
t417 cell_H25(.x1(D6), .y4(NET00190), .x5(CA), .x6(D14), .x10(CB));
t428 cell_K28(.x2(NET00148), .y3(NET00057));
t428 cell_K17(.x2(NET00249), .y3(NET00001));
t429 cell_K20(.y3(NET00007), .x5(NET00164));
t378 cell_L33(.x1(RC1), .y2(NET00199), .x3(NET00175), .x5(nRC0));
t429 cell_K32(.y3(NET00035), .x5(NET00146));
t416 cell_D39(.c1(NET00108), .q4(R1), .d5(D1));
t390 cell_M15(.x1(D10), .y4(NET00161), .x5(NET00165), .x6(D11), .y9(NET00233), .x10(NET00165));
t395 cell_G30(.x1(COM), .y2(NET00232), .x3(NET00232), .x4(NET00230), .x5(NET00230), .x6(COM), .y8(NET00170));
t416 cell_G39(.c1(NET00108), .q4(R3), .d5(D3));
t395 cell_I10(.x1(D7), .y2(NET00256), .x3(NET00256), .x4(NET00240), .x5(NET00240), .x6(D7), .y8(NET00209));
t395 cell_H30(.x1(COM), .y2(NET00222), .x3(NET00222), .x4(NET00220), .x5(NET00220), .x6(COM), .y8(NET00223));
t371 cell_H10(.x1(NET00129), .y3(nAD13), .y4(NET00128), .x6(NET00130));
t416 cell_I39(.c1(NET00108), .q4(R5), .d5(D5));
t395 cell_I12(.x1(D6), .y2(NET00257), .x3(NET00257), .x4(NET00239), .x5(NET00239), .x6(D6), .y8(NET00135));
t383 cell_H12(.x1(NET00132), .y2(NET00123), .x3(NET00133), .x4(NET00135), .x5(NET00131), .x6(NET00134));
t395 cell_G36(.x1(COM), .y2(NET00228), .x3(NET00228), .x4(NET00227), .x5(NET00227), .x6(COM), .y8(NET00229));
t416 cell_L39(.c1(NET00108), .q4(R7), .d5(D7));
t395 cell_I14(.x1(D5), .y2(NET00259), .x3(NET00259), .x4(NET00237), .x5(NET00237), .x6(D5), .y8(NET00134));
t395 cell_H36(.x1(COM), .y2(NET00226), .x3(NET00226), .x4(NET00224), .x5(NET00224), .x6(COM), .y8(NET00160));
t416 cell_N39(.c1(NET00035), .q4(R15), .d5(D15));
t378 cell_L24(.x1(RC1), .y2(NET00154), .x3(NET00155), .x5(nRC0));
t378 cell_L26(.x1(RC1), .y2(NET00152), .x3(NET00153), .x5(nRC0));
t378 cell_N28(.x1(NET00174), .y2(NET00156), .x3(nRC1), .x5(nRC0));
t378 cell_N26(.x1(NET00175), .y2(VIRQ), .x3(nRC1), .x5(nRC0));
t416 cell_M23(.c1(nCB), .q4(RIRQ), .d5(VIRQ));
t373 cell_J20(.x1(CA), .x3(CB), .y4(NET00164));
t374 cell_D9(.x1(NET00068), .x2(NET00067), .x3(nCD), .y4(PD1), .y8(NET00166));
t428 cell_E20(.x2(NET00203), .y3(NET00000));
t374 cell_D13(.x1(NET00074), .x2(NET00073), .x3(nCD), .y4(PD2), .y8(NET00186));
t395 cell_H18(.x1(COM), .y2(NET00121), .x3(NET00121), .x4(NET00119), .x5(NET00119), .x6(COM), .y8(NET00122));
t395 cell_G18(.x1(COM), .y2(NET00142), .x3(NET00142), .x4(NET00141), .x5(NET00141), .x6(COM), .y8(NET00143));
t395 cell_G8(.x1(D3), .y2(NET00171), .x3(NET00171), .x4(AD6), .x5(AD6), .x6(D3), .y8(NET00172));
t395 cell_G12(.x1(D1), .y2(NET00139), .x3(NET00139), .x4(AD4), .x5(AD4), .x6(D1), .y8(NET00133));
t395 cell_I8(.x1(D14), .y2(NET00236), .x3(NET00236), .x4(NET00214), .x5(NET00214), .x6(D14), .y8(NET00210));
t372 cell_J6(.x1(NET00252), .y2(NET00252), .y3(NET00253), .y4(NET00251), .x5(NET00251), .x6(NET00189));
t374 cell_I29(.x1(nRC0), .x2(RC3), .x3(nRC1), .y4(RC3), .y8(nRC3));
t390 cell_M13(.x1(D12), .y4(NET00235), .x5(NET00165), .x6(D13), .y9(NET00234), .x10(NET00165));
t429 cell_K9(.y3(nRC0), .x5(RC0));
t428 cell_K11(.x2(NET00250), .y3(RC1));
t428 cell_K24(.x2(NET00154), .y3(nCOM));
t384 cell_L23(.x1(NET00156), .y3(nDME3), .x5(RIRQ));
t380 cell_N24(.x1(NET00176), .y2(nCB), .y3(NET00260), .x4(nRC1), .x5(NET00260), .x6(nRC0));
t395 cell_H24(.x1(COM), .y2(NET00191), .x3(NET00191), .x4(NET00190), .x5(NET00190), .x6(COM), .y8(NET00192));
t395 cell_G24(.x1(COM), .y2(NET00195), .x3(NET00195), .x4(NET00194), .x5(NET00194), .x6(COM), .y8(NET00196));
t379 cell_L35(.x1(RC1), .y2(NET00167), .x3(NET00174), .y4(NET00198), .x5(nRC0), .x6(NET00174), .x8(RC0));
t372 cell_O31(.x1(NET00179), .y2(NET00179), .y3(NET00180), .y4(NET00178), .x5(NET00178), .x6(NET00181));
t429 cell_K25(.y3(COM), .x5(NET00154));
t428 cell_K31(.x2(NET00200), .y3(CB));
t428 cell_K27(.x2(NET00167), .y3(DME1));
t416 cell_M39(.c1(NET00035), .q4(R14), .d5(D14));
t416 cell_J39(.c1(NET00108), .q4(R6), .d5(D6));
t416 cell_H39(.c1(NET00108), .q4(R4), .d5(D4));
t416 cell_F39(.c1(NET00108), .q4(R2), .d5(D2));
t417 cell_H31(.x1(D5), .y4(NET00220), .x5(CA), .x6(D13), .x10(CB));
t417 cell_G31(.x1(D1), .y4(NET00230), .x5(CA), .x6(D9), .x10(CB));
t382 cell_H11(.x1(nAD13), .y2(NET00126), .x3(nRC3), .x4(NET00128), .x5(NET00123), .x6(NET00127), .y8(NET00127));
t417 cell_H37(.x1(D4), .y4(NET00224), .x5(CA), .x6(D12), .x10(CB));
t417 cell_G37(.x1(D0), .y4(NET00227), .x5(CA), .x6(D8), .x10(CB));
t372 cell_F20(.x1(NET00202), .y2(NET00202), .y3(NET00203), .y4(NET00201), .x5(NET00201), .x6(NET00204));
t416 cell_C39(.c1(NET00108), .q4(R0), .d5(D0));
t380 cell_N22(.x1(NET00153), .y2(nCA), .y3(NET00261), .x4(nRC1), .x5(NET00261), .x6(nRC0));
t378 cell_J19(.x1(NET00165), .y2(NET00246), .x3(NET00044), .x5(NET00007));
t383 cell_H9(.x1(NET00172), .y2(NET00130), .x3(NET00169), .x4(NET00211), .x5(NET00209), .x6(NET00210));
t374 cell_D5(.x1(NET00061), .x2(NET00060), .x3(nCD), .y4(PD0), .y8(NET00162));

endmodule
//______________________________________________________________________________
//
