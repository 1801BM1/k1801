//
// Copyright (c) 2013 by 1801BM1@gmail.com
//______________________________________________________________________________
//
`timescale 1ns / 100ps

module vp_128
(
   inout[15:0] PIN_nAD,       // Address/Data inverted bus
                              //
   input       PIN_nSYNC,     //
   input       PIN_nDIN,      //
   input       PIN_nDOUT,     //
   input       PIN_nINIT,     //
   input       PIN_CLK,       //
   output      PIN_nRPLY,     //
                              //
   output[3:0] PIN_nDS,       //
   output      PIN_nMSW,      //
   output      PIN_nST,       //
   output      PIN_DIR,       //
   output      PIN_HS,        //
   output      PIN_nWRE,      //
                              //
   output[3:1] PIN_nDO,       //
   output      PIN_nREZ,      //
   input       PIN_nDI,       //
   input       PIN_IND,       //
   input       PIN_TR0,       //
   input       PIN_RDY,       //
   input       PIN_WRP        //
);

//______________________________________________________________________________
//
// Autogenerated netlist
//
wire GND = 1'b0;
wire nBIT_CNT0;
wire nBIT_CNT2;
wire SREG4;
wire nSYNC;
wire CLK;
wire BCNT_CLK;
wire nAD1;
wire CRC_CLK0;
wire CRC_RST2;
wire CSR_TR;
wire nSTB_P09;
wire nLATCH_TR;
wire nSTB_P03;
wire SREG5;
wire WRE;
wire STB_P07;
wire OE_RDAT;
wire INIT_073;
wire MARKER;
wire DAT_WR_E4;
wire IND;
wire RDINIT0;
wire SREG6;
wire nSREG5;
wire nRDR_STB;
wire nDAT_RD;
wire nSREG7;
wire nRDR0;
wire nRDR9;
wire nAD15;
wire SREG_LD;
wire SEL_HB;
wire SREG_SH;
wire CRC_RST0;
wire nAD9;
wire nAD10;
wire nRDR13;
wire nRDR6;
wire nOE_RDAT;
wire nDAT_WR;
wire nRDR1;
wire SEL0;
wire nRDR2;
wire nRDR3;
wire CRC_CLK1;
wire nRDR4;
wire nCRC_CLK1;
wire nRDR5;
wire nAD2;
wire nCRC_RST;
wire CSR_WM;
wire CRC_IN0;
wire nSREG_Q;
wire nAD0;
wire nAD3;
wire nAD4;
wire nAD5;
wire nAD6;
wire nAD7;
wire nAD8;
wire nAD11;
wire nAD12;
wire nAD13;
wire nAD14;
wire SREG7;
wire nMARK_A1;
wire nWCLK;
wire nRDD_CLK;
wire STB_P11;
wire nAPC_CLK;
wire CRC_RST3;
wire OE_CSR;
wire INIT_F26;
wire PLL_RDY;
wire CRC_VALID;
wire nWCLK0;
wire nPLL_C;
wire APC_CLK;
wire SEL_LB;
wire SREG0;
wire PLL_EQ7;
wire nCLK;
wire PLL_S;
wire RDATA;
wire RDATA_Y;
wire nPLL_6OR7;
wire PLL_C;
wire nRDATA_Y;
wire STB_P15;
wire CRC_RST1;
wire DIN;
wire nRPLY;
wire nINIT;
wire RDINIT1;
wire WBIT2;
wire nCRC15;
wire PLL_H;
wire SREG_Q;
wire nRDR7;
wire nRDR8;
wire nRDR10;
wire nRDR11;
wire WRP;
wire nRDR12;
wire RDR_LSTB;
wire nRDR14;
wire nRDR15;
wire CSR_CRC;
wire RDR_HSTB;
wire nSREG_IN;
wire INIT_106;
wire nPLL_Z;
wire DOUT;
wire nSREG0;
wire SREG1;
wire SREG2;
wire SREG3;
wire SREG_SH_nLD;
wire nCRC_CLK0;
wire WBIT0;
wire LAST_WR;
wire nCSR_WR;
wire nCSR_RD;
wire PLL_CLK6;
wire PLL_A;
wire PLL_B;
wire PLL_2OR3;
wire nPLL_B;
wire SEL2;
wire RDR_STB;
wire nCSR_GDR;
wire CSR_GDR;
wire nPLL_A;
wire CRC15;
wire LATCH_TR;
wire FIN_STB;
wire RDD_CLK;
wire nWRE;
wire WBIT8;
wire nGDR;
wire MARK1;
wire MARK0;
wire STB_P09;
wire nWBIT0;
wire RDR_HSTB0;
wire WCLK;
wire RDR_LSTB0;
wire nWBIT1;
wire WBIT1;
wire MODE_R_nW;
wire WBIT3;
wire WBIT5;
wire WBIT4;
wire BIT_CNT0;
wire nBIT_CNT1;
wire MODE_nRn_W;
wire nSTB_P11;
wire PLL_B_DELAYED;
wire WBIT6;
wire PLL_B0;
wire nWBIT5;
wire nWBIT6;

wire NET00000;
wire NET00001;
wire NET00003;
wire NET00005;
wire NET00006;
wire NET00009;
wire NET00010;
wire NET00011;
wire NET00013;
wire NET00015;
wire NET00016;
wire NET00017;
wire NET00018;
wire NET00019;
wire NET00376;
wire NET00021;
wire NET00023;
wire NET00024;
wire NET00365;
wire NET00026;
wire NET00604;
wire NET00028;
wire NET00029;
wire NET00031;
wire NET00139;
wire NET00033;
wire NET00034;
wire NET00147;
wire NET00037;
wire NET00162;
wire NET00039;
wire NET00040;
wire NET00041;
wire NET00042;
wire NET00047;
wire NET00135;
wire NET00050;
wire NET00051;
wire NET00052;
wire NET00053;
wire NET00054;
wire NET00055;
wire NET00057;
wire NET00059;
wire NET00127;
wire NET00061;
wire NET00062;
wire NET00063;
wire NET00064;
wire NET00065;
wire NET00066;
wire NET00067;
wire NET00068;
wire NET00069;
wire NET00070;
wire NET00089;
wire NET00074;
wire NET00077;
wire NET00079;
wire NET00012;
wire NET00356;
wire NET00085;
wire NET00086;
wire NET00087;
wire NET00091;
wire NET00092;
wire NET00212;
wire NET00094;
wire NET00095;
wire NET00098;
wire NET00099;
wire NET00100;
wire NET00101;
wire NET00102;
wire NET00104;
wire NET00273;
wire NET00274;
wire NET00441;
wire NET00432;
wire NET00111;
wire NET00112;
wire NET00113;
wire NET00116;
wire NET00117;
wire NET00118;
wire NET00120;
wire NET00272;
wire NET00123;
wire NET00287;
wire NET00286;
wire NET00281;
wire NET00131;
wire NET00132;
wire NET00133;
wire NET00134;
wire NET00275;
wire NET00136;
wire NET00137;
wire NET00351;
wire NET00140;
wire NET00142;
wire NET00143;
wire NET00144;
wire NET00375;
wire NET00359;
wire NET00447;
wire NET00360;
wire NET00151;
wire NET00173;
wire NET00154;
wire NET00155;
wire NET00157;
wire NET00165;
wire NET00159;
wire NET00161;
wire NET00596;
wire NET00477;
wire NET00190;
wire NET00175;
wire NET00178;
wire NET00182;
wire NET00183;
wire NET00186;
wire NET00372;
wire NET00569;
wire NET00189;
wire NET00191;
wire NET00192;
wire NET00193;
wire NET00194;
wire NET00195;
wire NET00223;
wire NET00196;
wire NET00198;
wire NET00199;
wire NET00082;
wire NET00470;
wire NET00357;
wire NET00560;
wire NET00206;
wire NET00208;
wire NET00209;
wire NET00210;
wire NET00211;
wire NET00213;
wire NET00214;
wire NET00250;
wire NET00217;
wire NET00340;
wire NET00219;
wire NET00471;
wire NET00221;
wire NET00358;
wire NET00225;
wire NET00226;
wire NET00227;
wire NET00229;
wire NET00336;
wire NET00231;
wire NET00233;
wire NET00234;
wire NET00235;
wire NET00238;
wire NET00239;
wire NET00240;
wire NET00241;
wire NET00242;
wire NET00253;
wire NET00244;
wire NET00247;
wire NET00248;
wire NET00249;
wire NET00297;
wire NET00252;
wire NET00254;
wire NET00255;
wire NET00256;
wire NET00258;
wire NET00257;
wire NET00259;
wire NET00260;
wire NET00261;
wire NET00262;
wire NET00263;
wire NET00264;
wire NET00301;
wire NET00362;
wire NET00364;
wire NET00267;
wire NET00268;
wire NET00270;
wire NET00271;
wire NET00567;
wire NET00363;
wire NET00565;
wire NET00566;
wire NET00462;
wire NET00002;
wire NET00279;
wire NET00280;
wire NET00341;
wire NET00282;
wire NET00284;
wire NET00561;
wire NET00348;
wire NET00288;
wire NET00289;
wire NET00293;
wire NET00295;
wire NET00332;
wire NET00298;
wire NET00299;
wire NET00300;
wire NET00302;
wire NET00304;
wire NET00305;
wire NET00307;
wire NET00461;
wire NET00308;
wire NET00309;
wire NET00310;
wire NET00312;
wire NET00460;
wire NET00313;
wire NET00314;
wire NET00317;
wire NET00320;
wire NET00319;
wire NET00575;
wire NET00580;
wire NET00323;
wire NET00324;
wire NET00020;
wire NET00383;
wire NET00331;
wire NET00583;
wire NET00579;
wire NET00417;
wire NET00347;
wire NET00379;
wire NET00380;
wire NET00576;
wire NET00551;
wire NET00439;
wire NET00444;
wire NET00442;
wire NET00445;
wire NET00368;
wire NET00367;
wire NET00552;
wire NET00558;
wire NET00440;
wire NET00443;
wire NET00559;
wire NET00557;
wire NET00603;
wire NET00369;
wire NET00371;
wire NET00373;
wire NET00571;
wire NET00584;
wire NET00541;
wire NET00459;
wire NET00381;
wire NET00384;
wire NET00385;
wire NET00587;
wire NET00387;
wire NET00392;
wire NET00393;
wire NET00394;
wire NET00395;
wire NET00396;
wire NET00397;
wire NET00398;
wire NET00401;
wire NET00204;
wire NET00403;
wire NET00405;
wire NET00406;
wire NET00407;
wire NET00408;
wire NET00409;
wire NET00410;
wire NET00411;
wire NET00412;
wire NET00415;
wire NET00416;
wire NET00613;
wire NET00556;
wire NET00422;
wire NET00555;
wire NET00427;
wire NET00426;
wire NET00507;
wire NET00428;
wire NET00429;
wire NET00430;
wire NET00431;
wire NET00509;
wire NET00433;
wire NET00434;
wire NET00436;
wire NET00520;
wire NET00508;
wire NET00506;
wire NET00547;
wire NET00528;
wire NET00588;
wire NET00589;
wire NET00590;
wire NET00591;
wire NET00607;
wire NET00550;
wire NET00536;
wire NET00538;
wire NET00537;
wire NET00539;
wire NET00454;
wire NET00456;
wire NET00496;
wire NET00474;
wire NET00519;
wire NET00545;
wire NET00543;
wire NET00518;
wire NET00479;
wire NET00522;
wire NET00524;
wire NET00007;
wire NET00505;
wire NET00610;
wire NET00008;
wire NET00542;
wire NET00595;
wire NET00586;
wire NET00484;
wire NET00485;
wire NET00486;
wire NET00487;
wire NET00488;
wire NET00513;
wire NET00511;
wire NET00512;
wire NET00499;
wire NET00497;
wire NET00597;
wire NET00500;
wire NET00501;
wire NET00594;
wire NET00592;
wire NET00593;
wire NET00599;
wire NET00548;
wire NET00523;
wire NET00515;
wire NET00516;
wire NET00517;
wire NET00388;
wire NET00533;
wire NET00530;
wire NET00532;

//______________________________________________________________________________
//
// Autogenerated cell instantiations
//
tOUTPUT_OE  cell_PINOU1(.x1(NET00365),  .x2(NET00127), .y1(PIN_nAD[0]));
tOUTPUT_OE  cell_PINOU2(.x1(NET00147),  .x2(NET00127), .y1(PIN_nAD[1]));
tOUTPUT_OE  cell_PINOU3(.x1(NET00162),  .x2(NET00127), .y1(PIN_nAD[2]));
tOUTPUT_OE  cell_PINOU4(.x1(NET00165),  .x2(NET00135), .y1(PIN_nAD[3]));
tOUTPUT_OE  cell_PINOU5(.x1(NET00173),  .x2(NET00135), .y1(PIN_nAD[4]));
tOUTPUT_OE  cell_PINOU6(.x1(NET00360),  .x2(NET00135), .y1(PIN_nAD[5]));
tOUTPUT_OE  cell_PINOU7(.x1(NET00359),  .x2(NET00135), .y1(PIN_nAD[6]));
tOUTPUT_OE  cell_PINOU8(.x1(NET00356),  .x2(NET00127), .y1(PIN_nAD[7]));
tOUTPUT_OE  cell_PINOU9(.x1(NET00351),  .x2(NET00135), .y1(PIN_nAD[8]));
tOUTPUT_OE  cell_PINOU10(.x1(NET00275), .x2(NET00135), .y1(PIN_nAD[9]));
tOUTPUT_OE  cell_PINOU11(.x1(NET00281), .x2(NET00135), .y1(PIN_nAD[10]));
tOUTPUT_OE  cell_PINOU12(.x1(NET00286), .x2(NET00135), .y1(PIN_nAD[11]));
tOUTPUT_OE  cell_PINOU13(.x1(NET00287), .x2(NET00135), .y1(PIN_nAD[12]));
tOUTPUT_OE  cell_PINOU14(.x1(NET00272), .x2(NET00135), .y1(PIN_nAD[13]));
tOUTPUT_OE  cell_PINOU15(.x1(NET00273), .x2(NET00127), .y1(PIN_nAD[14]));
tOUTPUT_OE  cell_PINOU16(.x1(NET00274), .x2(NET00127), .y1(PIN_nAD[15]));

tINPUT      cell_PIN1(.y1(nAD0),   .x1(PIN_nAD[0]));
tINPUT      cell_PIN2(.y1(nAD1),   .x1(PIN_nAD[1]));
tINPUT      cell_PIN3(.y1(nAD2),   .x1(PIN_nAD[2]));
tINPUT      cell_PIN4(.y1(nAD3),   .x1(PIN_nAD[3]));
tINPUT      cell_PIN5(.y1(nAD4),   .x1(PIN_nAD[4]));
tINPUT      cell_PIN6(.y1(nAD5),   .x1(PIN_nAD[5]));
tINPUT      cell_PIN7(.y1(nAD6),   .x1(PIN_nAD[6]));
tINPUT      cell_PIN8(.y1(nAD7),   .x1(PIN_nAD[7]));
tINPUT      cell_PIN9(.y1(nAD8),   .x1(PIN_nAD[8]));
tINPUT      cell_PIN10(.y1(nAD9),  .x1(PIN_nAD[9]));
tINPUT      cell_PIN11(.y1(nAD10), .x1(PIN_nAD[10]));
tINPUT      cell_PIN12(.y1(nAD11), .x1(PIN_nAD[11]));
tINPUT      cell_PIN13(.y1(nAD12), .x1(PIN_nAD[12]));
tINPUT      cell_PIN14(.y1(nAD13), .x1(PIN_nAD[13]));
tINPUT      cell_PIN15(.y1(nAD14), .x1(PIN_nAD[14]));
tINPUT      cell_PIN16(.y1(nAD15), .x1(PIN_nAD[15]));

tINPUT      cell_PIN17(.y1(NET00444),  .x1(PIN_nSYNC));
tINPUT      cell_PIN18(.y1(NET00603),  .x1(PIN_nDIN));
tINPUT      cell_PIN19(.y1(NET00319),  .x1(PIN_nDOUT));
tINPUT      cell_PIN20(.y1(nINIT),     .x1(PIN_nINIT));
tINPUT      cell_PIN21(.y1(NET00376),  .x1(PIN_CLK));
tINPUT      cell_PIN24(.y1(IND),       .x1(PIN_IND));
tINPUT      cell_PIN29(.y2(NET00381),  .x1(PIN_nDI));
tINPUT      cell_PIN31(.y1(WRP),       .x1(PIN_WRP));
tINPUT      cell_PIN32(.y1(NET00139),  .x1(PIN_RDY));
tINPUT      cell_PIN33(.y1(NET00604),  .x1(PIN_TR0));

tOUTPUT_OC  cell_PIN23(.x1(nRPLY),     .y1(PIN_nRPLY));
tOUTPUT     cell_PIN25(.x1(NET00369),  .y1(PIN_nDO[3]));
tOUTPUT     cell_PIN26(.x1(NET00373),  .y1(PIN_nDO[2]));
tOUTPUT     cell_PIN27(.x1(NET00371),  .y1(PIN_nDO[1]));
tOUTPUT     cell_PIN28(.x1(nWRE),      .y1(PIN_nWRE));
tOUTPUT     cell_PIN30(.x1(NET00137),  .y1(PIN_nREZ));
tOUTPUT     cell_PIN34(.x1(NET00131),  .y1(PIN_nST));
tOUTPUT     cell_PIN35(.x1(NET00132),  .y1(PIN_DIR));
tOUTPUT     cell_PIN36(.x1(NET00133),  .y1(PIN_HS));
tOUTPUT     cell_PIN37(.x1(NET00136),  .y1(PIN_nMSW));
tOUTPUT     cell_PIN38(.x1(NET00143),  .y1(PIN_nDS[3]));
tOUTPUT     cell_PIN39(.x1(NET00144),  .y1(PIN_nDS[2]));
tOUTPUT     cell_PIN40(.x1(NET00257),  .y1(PIN_nDS[1]));
tOUTPUT     cell_PIN41(.x1(NET00575),  .y1(PIN_nDS[0]));

t387 cell_A35(.x1(WBIT8), .y2(NET00500), .x3(NET00532), .y4(NET00548), .x5(CSR_WM), .x6(NET00497));
t376 cell_A38(.x1(NET00548), .x3(NET00536), .y4(NET00369), .x6(NET00539), .x8(NET00537), .y9(NET00373));
t376 cell_B39(.x1(NET00501), .x3(NET00515), .y4(NET00536), .x6(NET00501), .x8(NET00516), .y9(NET00537));
t406 cell_L34(.c1(CRC_CLK1), .r2(CRC_RST3), .q3(NET00304), .q4(NET00301), .r5(NET00310), .s10(NET00308));
t416 cell_A0(.c1(RDR_HSTB), .q4(NET00272), .d5(nRDR13));
t417 cell_A1(.x1(CSR_CRC), .y4(NET00273), .x5(NET00140), .x6(NET00432), .x10(OE_RDAT));
t429 cell_K3(.y3(NET00127), .x5(OE_CSR));
t388 cell_A10(.x1(DOUT), .y2(NET00317), .x3(DIN), .y4(NET00267), .y5(NET00314), .x6(DOUT), .x7(NET00314), .x10(nRPLY));
t376 cell_A11(.x1(nSYNC), .x3(NET00603), .y4(DIN), .x6(nSYNC), .x8(NET00319), .y9(DOUT));
t373 cell_H36(.x1(NET00396), .x3(NET00408), .y4(NET00410));
t370 cell_B27(.y2(NET00416), .x5(nSTB_P03));
t377 cell_A23(.x1(nPLL_6OR7), .y2(NET00426), .x3(nPLL_A), .y4(PLL_EQ7), .x5(nPLL_A), .x6(nPLL_6OR7), .x8(NET00403), .y9(PLL_CLK6));
t379 cell_A26(.x1(NET00428), .y2(NET00430), .x3(NET00429), .y4(NET00428), .x5(PLL_S), .x6(NET00430), .x8(NET00206));
t406 cell_G32(.c1(RDATA), .r2(RDD_CLK), .q4(nSREG_IN), .r5(GND), .s10(nRDD_CLK));
t379 cell_D24(.x1(NET00393), .y2(NET00395), .x3(PLL_B), .y4(NET00393), .x5(NET00392), .x6(NET00395), .x8(nPLL_C));
t406 cell_G24(.c1(STB_P15), .r2(INIT_106), .q3(NET00217), .q4(NET00249), .r5(NET00288), .s10(NET00289));
t376 cell_G23(.x1(NET00298), .x3(NET00299), .y4(NET00300), .x6(NET00300), .x8(NET00002), .y9(NET00299));
t429 cell_E37(.y3(NET00474), .x5(nWCLK));
t428 cell_E35(.x2(NET00376), .y3(CLK));
t429 cell_E36(.y3(nWCLK0), .x5(WCLK));
t376 cell_C2(.x1(SREG7), .x3(NET00094), .y4(nRDR15), .x6(SREG7), .x8(NET00095), .y9(nRDR7));
t416 cell_B1(.c1(RDR_HSTB), .q3(NET00432), .d5(nRDR14));
t416 cell_B2(.c1(RDR_HSTB), .q3(NET00441), .d5(nRDR15));
t416 cell_L5(.c1(NET00477), .q3(NET00116), .d5(nAD4));
t390 cell_L4(.x1(nAD2), .y4(NET00367), .x5(nAD5), .x6(nAD7), .y9(NET00368), .x10(nAD8));
t374 cell_B10(.x1(NET00270), .x2(NET00267), .x3(NET00267), .y4(NET00268), .y8(NET00271));
t406 cell_B11(.c1(CLK), .r2(NET00267), .q4(nRPLY), .r5(GND), .s10(NET00268));
t377 cell_B18(.x1(nRDATA_Y), .y2(PLL_2OR3), .x3(PLL_2OR3), .y4(NET00284), .x5(NET00282), .x6(NET00284), .x8(PLL_H), .y9(NET00204));
t387 cell_I39(.x1(NET00397), .y2(nCRC_RST), .x3(NET00398), .y4(NET00396), .x5(NET00396), .x6(FIN_STB));
t390 cell_D31(.x1(MARK0), .y4(nMARK_A1), .x5(MARK1), .x6(WRE), .y9(nWCLK), .x10(NET00416));
t428 cell_E18(.x2(SEL_LB), .y3(NET00099));
t377 cell_F26(.x1(INIT_F26), .y2(INIT_F26), .x3(NET00293), .y4(NET00331), .x5(nINIT), .x6(NET00295), .x8(NET00002), .y9(NET00293));
t379 cell_A24(.x1(NET00429), .y2(NET00431), .x3(NET00206), .y4(NET00429), .x5(NET00428), .x6(NET00431), .x8(NET00426));
t413 cell_L23(.q1(LAST_WR), .r3(INIT_073), .q4(NET00020), .r5(nOE_RDAT), .x7(DAT_WR_E4), .y8(NET00074), .s10(NET00074));
t374 cell_B30(.x1(PLL_RDY), .x2(RDR_STB), .x3(MODE_nRn_W), .y4(NET00244), .y8(nRDR_STB));
t428 cell_E33(.x2(NET00479), .y3(MODE_nRn_W));
t406 cell_B37(.c1(NET00474), .r2(nWRE), .q3(WBIT5), .q4(nWBIT5), .r5(NET00519), .s10(WBIT4));
t406 cell_B36(.c1(nWCLK0), .r2(nWRE), .q3(WBIT6), .q4(nWBIT6), .r5(nWBIT5), .s10(WBIT5));
t406 cell_D37(.c1(NET00474), .r2(nWRE), .q3(WBIT1), .q4(nWBIT1), .r5(nWBIT0), .s10(WBIT0));
t416 cell_F0(.c1(RDR_HSTB), .q4(NET00281), .d5(nRDR10));
t376 cell_F2(.x1(SREG5), .x3(NET00094), .y4(nRDR13), .x6(SREG5), .x8(NET00095), .y9(nRDR5));
t376 cell_D2(.x1(SREG6), .x3(NET00094), .y4(nRDR14), .x6(SREG6), .x8(NET00095), .y9(nRDR6));
t416 cell_M5(.c1(NET00477), .q3(NET00357), .d5(nAD3));
t416 cell_M4(.c1(NET00477), .q3(NET00470), .d5(nAD2));
t406 cell_C12(.c1(NET00011), .r2(INIT_073), .q3(SREG_Q), .q4(nSREG_Q), .r5(nSREG7), .s10(SREG7));
t408 cell_M12(.q2(CSR_TR), .r5(NET00513), .s10(NET00511));
t376 cell_A28(.x1(NET00436), .x3(NET00077), .y4(NET00433), .x6(RDINIT0), .x8(NET00433), .y9(NET00436));
t428 cell_E19(.x2(SEL_LB), .y3(NET00095));
t379 cell_I19(.x1(nBIT_CNT0), .y2(BIT_CNT0), .x3(NET00212), .y4(nBIT_CNT0), .x5(RDINIT1), .x6(BIT_CNT0), .x8(NET00583));
t379 cell_H19(.x1(nBIT_CNT1), .y2(NET00599), .x3(NET00000), .y4(nBIT_CNT1), .x5(RDINIT1), .x6(NET00599), .x8(NET00003));
t379 cell_A30(.x1(NET00542), .y2(PLL_RDY), .x3(NET00433), .y4(NET00542), .x5(RDINIT0), .x6(PLL_RDY), .x8(NET00434));
t406 cell_F25(.c1(RDATA), .r2(nRDD_CLK), .q3(NET00289), .q4(NET00288), .r5(GND), .s10(RDD_CLK));
t428 cell_E23(.x2(NET00299), .y3(PLL_H));
t416 cell_A7(.c1(NET00442), .q3(SEL2), .q4(SEL0), .d5(nAD1));
t428 cell_E38(.x2(NET00456), .y3(nWRE));
t376 cell_A39(.x1(NET00538), .x3(NET00550), .y4(NET00371), .x6(NET00501), .x8(NET00517), .y9(NET00550));
t429 cell_E39(.y3(NET00219), .x5(nCSR_WR));
t416 cell_I0(.c1(RDR_HSTB), .q4(NET00351), .d5(nRDR8));
t376 cell_H2(.x1(SREG3), .x3(NET00094), .y4(nRDR11), .x6(SREG3), .x8(NET00095), .y9(nRDR3));
t416 cell_N4(.c1(NET00477), .q3(NET00372), .d5(nAD0));
t380 cell_N3(.x1(nAD6), .y2(NET00558), .y3(NET00576), .x4(nAD4), .x5(NET00576), .x6(nAD3));
t406 cell_D12(.c1(NET00011), .r2(INIT_073), .q4(NET00111), .r5(NET00199), .s10(SREG6));
t379 cell_O19(.x1(NET00485), .y2(NET00488), .x3(NET00487), .y4(NET00485), .x5(FIN_STB), .x6(NET00488), .x8(RDR_HSTB));
t428 cell_K18(.x2(NET00484), .y3(nLATCH_TR));
t379 cell_G19(.x1(nBIT_CNT2), .y2(NET00597), .x3(NET00053), .y4(nBIT_CNT2), .x5(RDINIT1), .x6(NET00597), .x8(NET00055));
t379 cell_F19(.x1(SEL_LB), .y2(SEL_HB), .x3(NET00089), .y4(SEL_LB), .x5(RDINIT1), .x6(SEL_HB), .x8(NET00091));
t379 cell_F18(.x1(NET00092), .y2(NET00091), .x3(NET00597), .y4(NET00092), .x5(NET00089), .x6(NET00091), .x8(SEL_LB));
t406 cell_H22(.c1(STB_P15), .r2(INIT_106), .q3(NET00210), .q4(NET00208), .r5(NET00247), .s10(NET00248));
t387 cell_H25(.x1(NET00020), .y2(NET00252), .x3(nMARK_A1), .y4(MARKER), .x5(NET00012), .x6(NET00252));
t376 cell_C39(.x1(NET00506), .x3(NET00007), .y4(NET00520), .x6(NET00381), .x8(NET00520), .y9(NET00506));
t429 cell_K0(.y3(NET00135), .x5(OE_RDAT));
t429 cell_K2(.y3(OE_RDAT), .x5(nDAT_RD));
t384 cell_J2(.x1(nDAT_RD), .y3(OE_CSR), .x5(nCSR_RD));
t417 cell_O3(.x1(WRP), .y4(NET00162), .x5(NET00140), .x6(NET00157), .x10(OE_RDAT));
t416 cell_O4(.c1(RDR_LSTB), .q3(NET00157), .d5(nRDR2));
t418 cell_F9(.x1(NET00050), .x2(NET00087), .y3(NET00086), .y4(NET00087), .x5(SREG_SH), .x6(NET00561), .x10(SREG_LD));
t379 cell_I18(.x1(NET00213), .y2(NET00583), .x3(BCNT_CLK), .y4(NET00213), .x5(NET00212), .x6(NET00583), .x8(nBIT_CNT0));
t379 cell_I20(.x1(NET00212), .y2(NET00214), .x3(NET00213), .y4(NET00212), .x5(RDINIT1), .x6(NET00214), .x8(BCNT_CLK));
t379 cell_N22(.x1(MODE_R_nW), .y2(NET00479), .x3(NET00592), .y4(MODE_R_nW), .x5(INIT_073), .x6(NET00479), .x8(NET00594));
t379 cell_H18(.x1(NET00001), .y2(NET00003), .x3(BIT_CNT0), .y4(NET00001), .x5(NET00000), .x6(NET00003), .x8(nBIT_CNT1));
t406 cell_I22(.c1(STB_P15), .r2(INIT_106), .q3(NET00161), .q4(NET00159), .r5(NET00211), .s10(NET00209));
t429 cell_E30(.y3(STB_P07), .x5(NET00412));
t429 cell_E26(.y3(PLL_S), .x5(NET00331));
t406 cell_D36(.c1(nWCLK0), .r2(nWRE), .q3(WBIT2), .q4(NET00496), .r5(nWBIT1), .s10(WBIT1));
t406 cell_L28(.c1(CRC_CLK1), .r2(CRC_RST3), .q3(NET00059), .q4(NET00062), .r5(NET00057), .s10(NET00061));
t416 cell_M0(.c1(RDR_LSTB), .q4(NET00359), .d5(nRDR6));
t417 cell_L0(.x1(CSR_TR), .y4(NET00356), .x5(NET00140), .x6(NET00375), .x10(OE_RDAT));
t376 cell_L2(.x1(SREG1), .x3(NET00094), .y4(nRDR9), .x6(SREG1), .x8(NET00095), .y9(nRDR1));
t371 cell_A6(.x1(NET00444), .y3(NET00447), .y4(NET00442), .x6(NET00447));
t418 cell_H9(.x1(NET00347), .x2(NET00009), .y3(NET00005), .y4(NET00009), .x5(SREG_SH), .x6(NET00348), .x10(SREG_LD));
t379 cell_H20(.x1(NET00000), .y2(NET00250), .x3(NET00001), .y4(NET00000), .x5(RDINIT1), .x6(NET00250), .x8(BIT_CNT0));
t385 cell_D19(.x1(NET00204), .x2(CLK), .y3(NET00206), .x5(CLK), .y8(nCLK));
t429 cell_E24(.y3(STB_P15), .x5(NET00280));
t379 cell_A18(.x1(NET00324), .y2(NET00610), .x3(nPLL_Z), .y4(NET00324), .x5(NET00323), .x6(NET00610), .x8(APC_CLK));
t379 cell_A19(.x1(APC_CLK), .y2(nAPC_CLK), .x3(NET00323), .y4(APC_CLK), .x5(RDINIT0), .x6(nAPC_CLK), .x8(NET00610));
t406 cell_J22(.c1(STB_P15), .r2(INIT_106), .q4(NET00155), .r5(NET00151), .s10(NET00154));
t378 cell_C24(.x1(PLL_H), .y2(nPLL_B), .x3(NET00406), .x5(PLL_B));
t381 cell_F23(.x1(PLL_B_DELAYED), .y2(NET00298), .x3(PLL_C), .x4(NET00293), .x6(nRDATA_Y));
t376 cell_B38(.x1(NET00497), .x3(NET00533), .y4(NET00538), .x6(NET00497), .x8(NET00530), .y9(NET00539));
t418 cell_D32(.x1(nLATCH_TR), .x2(WBIT0), .y3(nWBIT0), .y4(WBIT0), .x5(nSREG_Q), .x6(CRC15), .x10(LATCH_TR));
t379 cell_D39(.x1(NET00506), .y2(NET00508), .x3(NET00507), .y4(NET00507), .x5(NET00381), .x6(NET00508), .x8(CLK));
t416 cell_O0(.c1(RDR_LSTB), .q4(NET00173), .d5(nRDR4));
t416 cell_N0(.c1(RDR_LSTB), .q4(NET00360), .d5(nRDR5));
t379 cell_B6(.x1(NET00556), .y2(NET00555), .x3(CLK), .y4(NET00556), .x5(NET00613), .x6(NET00555), .x8(NET00271));
t418 cell_J9(.x1(NET00541), .x2(NET00566), .y3(NET00565), .y4(NET00566), .x5(SREG_SH), .x6(NET00567), .x10(SREG_LD));
t379 cell_G18(.x1(NET00054), .y2(NET00055), .x3(NET00599), .y4(NET00054), .x5(NET00053), .x6(NET00055), .x8(nBIT_CNT2));
t371 cell_F24(.x1(NET00279), .y3(nRDD_CLK), .y4(RDD_CLK), .x6(nRDD_CLK));
t377 cell_C18(.x1(nSTB_P09), .y2(nSTB_P09), .x3(NET00244), .y4(BCNT_CLK), .x5(STB_P09), .x6(PLL_C), .x8(nAPC_CLK), .y9(STB_P09));
t379 cell_D26(.x1(NET00392), .y2(NET00394), .x3(NET00393), .y4(NET00392), .x5(PLL_S), .x6(NET00394), .x8(PLL_B));
t406 cell_N36(.c1(CRC_CLK1), .r2(CRC_RST1), .q3(NET00070), .q4(NET00069), .r5(NET00231), .s10(NET00229));
t428 cell_K23(.x2(INIT_106), .y3(INIT_073));
t380 cell_A34(.x1(CSR_WM), .y2(NET00532), .y3(NET00547), .x4(WBIT6), .x5(NET00547), .x6(nWBIT0));
t391 cell_M15(.x1(RDR_HSTB0), .x2(RDINIT0), .y3(NET00522), .y4(NET00523), .x5(LATCH_TR), .x6(NET00522), .y9(NET00524), .x10(NET00523));
t391 cell_D30(.x1(RDR_STB), .x2(nMARK_A1), .y3(NET00505), .y4(SREG_SH_nLD), .x5(MODE_nRn_W), .x6(RDR_STB), .y9(NET00398), .x10(NET00505));
t406 cell_C37(.c1(NET00474), .r2(nWRE), .q3(WBIT3), .q4(NET00518), .r5(NET00496), .s10(WBIT2));
t418 cell_D9(.x1(NET00085), .x2(NET00198), .y3(NET00196), .y4(NET00198), .x5(SREG_SH), .x6(NET00341), .x10(SREG_LD));
t416 cell_O1(.c1(RDR_LSTB), .q4(NET00165), .d5(nRDR3));
t429 cell_E7(.y3(SREG_LD), .x5(SREG_SH_nLD));
t429 cell_E12(.y3(NET00006), .x5(NET00134));
t373 cell_A29(.x1(NET00077), .x3(NET00433), .y4(NET00434));
t379 cell_A25(.x1(PLL_A), .y2(nPLL_A), .x3(NET00428), .y4(PLL_A), .x5(PLL_S), .x6(nPLL_A), .x8(NET00431));
t381 cell_G15(.x1(LATCH_TR), .y2(NET00017), .x3(nBIT_CNT1), .x4(nSTB_P11), .x6(BIT_CNT0));
t386 cell_F38(.x1(NET00454), .y2(NET00454), .y3(WRE), .y4(NET00456), .x5(MODE_nRn_W), .x6(WRP), .x7(NET00456));
t371 cell_F35(.x1(NET00007), .y3(NET00008), .y4(RDATA), .x6(NET00008));
t417 cell_C7(.x1(NET00099), .y4(NET00102), .x5(NET00098), .x6(NET00101), .x10(NET00100));
t428 cell_K12(.x2(STB_P15), .y3(NET00011));
t406 cell_H11(.c1(NET00006), .r2(NET00082), .q3(SREG3), .q4(NET00010), .r5(NET00005), .s10(NET00009));
t387 cell_N15(.x1(RDR_LSTB0), .y2(NET00511), .x3(RDINIT0), .y4(NET00513), .x5(nLATCH_TR), .x6(NET00512));
t418 cell_B12(.x1(STB_P07), .x2(nSTB_P11), .y3(STB_P11), .y4(NET00134), .x5(SREG_SH), .x6(STB_P11), .x10(SREG_LD));
t379 cell_O17(.x1(NET00487), .y2(NET00486), .x3(RDR_HSTB), .y4(NET00487), .x5(NET00485), .x6(NET00486), .x8(CSR_TR));
t379 cell_O18(.x1(NET00484), .y2(LATCH_TR), .x3(NET00485), .y4(NET00484), .x5(FIN_STB), .x6(LATCH_TR), .x8(NET00486));
t406 cell_F39(.c1(NET00219), .r2(NET00182), .q4(NET00137), .r5(nAD10), .s10(NET00379));
t416 cell_O10(.c1(RDR_LSTB), .q3(NET00142), .d5(nRDR0));
t418 cell_L9(.x1(nSREG_IN), .x2(NET00363), .y3(NET00362), .y4(NET00363), .x5(SREG_SH), .x6(NET00364), .x10(SREG_LD));
t382 cell_B3(.x1(nAD9), .y2(NET00551), .x3(nAD11), .x4(nAD10), .x5(NET00551), .x6(nAD12), .y8(NET00552));
t379 cell_B9(.x1(NET00270), .y2(NET00559), .x3(NET00613), .y4(NET00270), .x5(nSYNC), .x6(NET00559), .x8(NET00555));
t380 cell_A3(.x1(nAD15), .y2(NET00440), .y3(NET00439), .x4(nAD14), .x5(NET00439), .x6(nAD13));
t379 cell_B7(.x1(NET00613), .y2(NET00557), .x3(NET00556), .y4(NET00613), .x5(nSYNC), .x6(NET00557), .x8(CLK));
t428 cell_K15(.x2(NET00524), .y3(FIN_STB));
t394 cell_G26(.x1(RDATA_Y), .y2(NET00002), .x3(NET00293), .y4(NET00295), .x5(PLL_EQ7), .x6(PLL_EQ7), .y9(nPLL_Z), .x10(RDATA_Y));
t380 cell_B33(.x1(nWBIT6), .y2(NET00530), .y3(NET00528), .x4(WBIT0), .x5(NET00528), .x6(CSR_WM));
t383 cell_B4(.x1(NET00440), .y2(NET00445), .x3(NET00558), .x4(NET00552), .x5(NET00368), .x6(NET00367));
t384 cell_A4(.x1(NET00443), .y3(nSYNC), .x5(NET00447));
t390 cell_A9(.x1(SEL0), .y4(nCSR_WR), .x5(NET00317), .x6(SEL0), .y9(nCSR_RD), .x10(DIN));
t418 cell_O11(.x1(NET00604), .x2(OE_RDAT), .y3(nOE_RDAT), .y4(NET00365), .x5(NET00140), .x6(NET00142), .x10(OE_RDAT));
t406 cell_C36(.c1(nWCLK0), .r2(nWRE), .q3(WBIT4), .q4(NET00519), .r5(NET00518), .s10(WBIT3));
t416 cell_D5(.c1(DAT_WR_E4), .q3(NET00117), .d5(nAD12));
t416 cell_D4(.c1(DAT_WR_E4), .q3(NET00336), .d5(nAD13));
t381 cell_I5(.x1(SREG3), .y2(MARK0), .x3(SREG2), .x4(nSREG0), .x6(SREG1));
t429 cell_E4(.y3(DAT_WR_E4), .x5(nDAT_WR));
t406 cell_N30(.c1(CRC_CLK0), .r2(CRC_RST2), .q3(NET00225), .q4(NET00192), .r5(NET00235), .s10(NET00233));
t390 cell_C35(.x1(WBIT5), .y4(NET00515), .x5(nWBIT1), .x6(NET00516), .y9(NET00517), .x10(NET00515));
t406 cell_N26(.c1(CRC_CLK0), .r2(CRC_RST0), .q3(NET00589), .q4(NET00241), .r5(NET00590), .s10(NET00591));
t416 cell_O6(.c1(RDR_LSTB), .q3(NET00596), .d5(nRDR1));
t416 cell_G4(.c1(DAT_WR_E4), .q3(NET00123), .d5(nAD9));
t406 cell_A37(.c1(NET00474), .r2(nWRE), .q3(NET00545), .q4(NET00543), .r5(nWBIT6), .s10(WBIT6));
t406 cell_M36(.c1(CRC_CLK1), .r2(CRC_RST1), .q3(NET00607), .q4(NET00240), .r5(NET00256), .s10(NET00258));
t406 cell_A36(.c1(nWCLK0), .r2(nWRE), .q3(WBIT8), .r5(NET00543), .s10(NET00545));
t416 cell_G5(.c1(DAT_WR_E4), .q3(NET00120), .d5(nAD8));
t417 cell_L7(.x1(NET00099), .y4(NET00364), .x5(NET00372), .x6(NET00101), .x10(NET00120));
t406 cell_M34(.c1(CRC_CLK1), .r2(CRC_RST1), .q3(NET00255), .q4(NET00242), .r5(NET00259), .s10(NET00260));
t406 cell_M28(.c1(CRC_CLK0), .r2(CRC_RST2), .q3(NET00026), .q4(NET00028), .r5(NET00024), .s10(NET00021));
t417 cell_I7(.x1(NET00099), .y4(NET00462), .x5(NET00470), .x6(NET00101), .x10(NET00471));
t416 cell_H5(.c1(NET00477), .q3(NET00340), .d5(nAD6));
t406 cell_M22(.c1(CRC_CLK0), .r2(CRC_RST0), .q3(NET00033), .q4(NET00029), .r5(NET00041), .s10(NET00039));
t429 cell_K27(.y3(CRC_RST0), .x5(nCRC_RST));
t406 cell_I11(.c1(NET00006), .r2(NET00082), .q3(SREG2), .q4(NET00584), .r5(NET00460), .s10(NET00461));
t417 cell_H7(.x1(NET00099), .y4(NET00348), .x5(NET00357), .x6(NET00101), .x10(NET00358));
t406 cell_F12(.c1(NET00011), .r2(INIT_073), .q4(NET00085), .r5(nSREG5), .s10(SREG5));
t406 cell_O27(.c1(NET00175), .r2(NET00182), .q4(NET00257), .r5(nAD1), .s10(NET00579));
t372 cell_O26(.x1(nAD2), .y2(NET00580), .y3(NET00189), .y4(NET00579), .x5(nAD0), .x6(nAD1));
t406 cell_J11(.c1(NET00006), .r2(NET00082), .q3(SREG1), .q4(NET00571), .r5(NET00565), .s10(NET00566));
t417 cell_F7(.x1(NET00099), .y4(NET00561), .x5(NET00560), .x6(NET00101), .x10(NET00336));
t417 cell_G7(.x1(NET00099), .y4(NET00118), .x5(NET00116), .x6(NET00101), .x10(NET00117));
t378 cell_C25(.x1(nPLL_B), .y2(PLL_B), .x3(NET00405), .x5(PLL_S));
t379 cell_A20(.x1(NET00323), .y2(NET00427), .x3(NET00324), .y4(NET00323), .x5(RDINIT0), .x6(NET00427), .x8(nPLL_Z));
t376 cell_I2(.x1(SREG2), .x3(NET00094), .y4(nRDR10), .x6(SREG2), .x8(NET00095), .y9(nRDR2));
t416 cell_J0(.c1(RDR_LSTB), .q3(NET00375), .d5(nRDR7));
t416 cell_H0(.c1(RDR_HSTB), .q4(NET00275), .d5(nRDR9));
t416 cell_D0(.c1(RDR_HSTB), .q4(NET00286), .d5(nRDR11));
t416 cell_B0(.c1(RDR_HSTB), .q4(NET00287), .d5(nRDR12));
t376 cell_G2(.x1(SREG4), .x3(NET00094), .y4(nRDR12), .x6(SREG4), .x8(NET00095), .y9(nRDR4));
t417 cell_A2(.x1(IND), .y4(NET00274), .x5(NET00140), .x6(NET00441), .x10(OE_RDAT));
t429 cell_K4(.y3(NET00140), .x5(nCSR_RD));
t406 cell_C11(.c1(NET00006), .r2(INIT_073), .q3(SREG7), .q4(nSREG7), .r5(NET00112), .s10(NET00113));
t428 cell_E9(.x2(SREG_SH_nLD), .y3(SREG_SH));
t406 cell_D11(.c1(NET00006), .r2(INIT_073), .q3(SREG6), .q4(NET00199), .r5(NET00196), .s10(NET00198));
t376 cell_L15(.x1(nRDR_STB), .x3(NET00095), .y4(RDR_LSTB0), .x6(nRDR_STB), .x8(NET00094), .y9(RDR_HSTB0));
t428 cell_E20(.x2(SEL_HB), .y3(NET00094));
t387 cell_I15(.x1(BCNT_CLK), .y2(NET00586), .x3(NET00016), .y4(RDR_STB), .x5(nBIT_CNT0), .x6(NET00586));
t428 cell_E17(.x2(SEL_HB), .y3(NET00101));
t376 cell_G37(.x1(NET00422), .x3(NET00396), .y4(NET00408), .x6(FIN_STB), .x8(NET00408), .y9(NET00422));
t406 cell_H23(.c1(STB_P07), .r2(INIT_106), .q3(NET00248), .q4(NET00247), .r5(NET00249), .s10(NET00217));
t379 cell_N21(.x1(NET00593), .y2(NET00594), .x3(NET00018), .y4(NET00593), .x5(NET00592), .x6(NET00594), .x8(LAST_WR));
t391 cell_B20(.x1(PLL_2OR3), .x2(APC_CLK), .y3(NET00411), .y4(nSTB_P03), .x5(NET00411), .x6(PLL_CLK6), .y9(NET00412), .x10(NET00411));
t381 cell_I25(.x1(NET00155), .y2(NET00012), .x3(NET00161), .x4(NET00217), .x6(NET00208));
t429 cell_E27(.y3(INIT_106), .x5(nINIT));
t390 cell_D33(.x1(nWCLK0), .y4(NET00501), .x5(WBIT3), .x6(WRE), .y9(WCLK), .x10(STB_P11));
t418 cell_C9(.x1(NET00111), .x2(NET00113), .y3(NET00112), .y4(NET00113), .x5(SREG_SH), .x6(NET00102), .x10(SREG_LD));
t417 cell_D7(.x1(NET00099), .y4(NET00341), .x5(NET00340), .x6(NET00101), .x10(NET00104));
t416 cell_J4(.c1(NET00477), .q3(NET00560), .d5(nAD5));
t376 cell_M2(.x1(SREG0), .x3(NET00094), .y4(nRDR8), .x6(SREG0), .x8(NET00095), .y9(nRDR0));
t429 cell_K37(.y3(CRC_RST1), .x5(nCRC_RST));
t406 cell_L11(.c1(NET00006), .r2(NET00082), .q3(SREG0), .q4(nSREG0), .r5(NET00362), .s10(NET00363));
t406 cell_G11(.c1(NET00006), .r2(NET00082), .q3(SREG4), .q4(NET00047), .r5(NET00051), .s10(NET00052));
t390 cell_A8(.x1(SEL2), .y4(nDAT_RD), .x5(DIN), .x6(SEL2), .y9(nDAT_WR), .x10(NET00317));
t418 cell_I9(.x1(NET00459), .x2(NET00461), .y3(NET00460), .y4(NET00461), .x5(SREG_SH), .x6(NET00462), .x10(SREG_LD));
t418 cell_G9(.x1(NET00013), .x2(NET00052), .y3(NET00051), .y4(NET00052), .x5(SREG_SH), .x6(NET00118), .x10(SREG_LD));
t381 cell_D13(.x1(nSREG7), .y2(MARK1), .x3(SREG4), .x4(SREG6), .x6(nSREG5));
t387 cell_A12(.x1(DOUT), .y2(NET00131), .x3(SEL2), .y4(NET00320), .x5(NET00320), .x6(nAD7));
t374 cell_M21(.x1(NET00042), .x2(IND), .x3(STB_P09), .y4(NET00015), .y8(NET00042));
t379 cell_G20(.x1(NET00053), .y2(NET00297), .x3(NET00054), .y4(NET00053), .x5(RDINIT1), .x6(NET00297), .x8(NET00599));
t379 cell_F20(.x1(NET00089), .y2(NET00332), .x3(NET00092), .y4(NET00089), .x5(RDINIT1), .x6(NET00332), .x8(NET00597));
t391 cell_B19(.x1(NET00279), .x2(nAPC_CLK), .y3(NET00279), .y4(nSTB_P11), .x5(PLL_2OR3), .x6(NET00279), .y9(NET00280), .x10(PLL_CLK6));
t378 cell_B25(.x1(PLL_H), .y2(NET00405), .x3(PLL_A), .x5(NET00415));
t379 cell_D25(.x1(nPLL_C), .y2(PLL_C), .x3(NET00392), .y4(nPLL_C), .x5(PLL_S), .x6(PLL_C), .x8(NET00395));
t406 cell_I23(.c1(STB_P07), .r2(INIT_106), .q3(NET00209), .q4(NET00211), .r5(NET00208), .s10(NET00210));
t406 cell_O23(.c1(NET00175), .r2(NET00182), .q4(NET00575), .r5(nAD0), .s10(NET00580));
t406 cell_J23(.c1(STB_P07), .r2(INIT_106), .q3(NET00154), .q4(NET00151), .r5(NET00159), .s10(NET00161));
t417 cell_J36(.x1(MODE_R_nW), .y4(CSR_CRC), .x5(NET00388), .x6(nLATCH_TR), .x10(MODE_nRn_W));
t429 cell_K35(.y3(CRC_RST2), .x5(nCRC_RST));
t418 cell_G27(.x1(nCLK), .x2(RDATA_Y), .y3(nRDATA_Y), .y4(RDATA_Y), .x5(NET00008), .x6(NET00008), .x10(nRDATA_Y));
t390 cell_B35(.x1(nWBIT5), .y4(NET00516), .x5(WBIT1), .x6(NET00532), .y9(NET00533), .x10(NET00530));
t379 cell_D38(.x1(NET00381), .y2(NET00007), .x3(NET00509), .y4(NET00509), .x5(CLK), .x6(NET00007), .x8(NET00508));
t406 cell_L12(.c1(STB_P15), .r2(NET00082), .q4(NET00541), .r5(nSREG0), .s10(SREG0));
t428 cell_K13(.x2(RDR_LSTB0), .y3(RDR_LSTB));
t406 cell_H12(.c1(NET00011), .r2(NET00082), .q4(NET00013), .r5(NET00010), .s10(SREG3));
t428 cell_E11(.x2(INIT_073), .y3(NET00082));
t428 cell_K19(.x2(RDR_HSTB0), .y3(RDR_HSTB));
t416 cell_C5(.c1(DAT_WR_E4), .q3(NET00104), .d5(nAD14));
t416 cell_C4(.c1(DAT_WR_E4), .q3(NET00100), .d5(nAD15));
t416 cell_N5(.c1(NET00477), .q3(NET00569), .d5(nAD1));
t416 cell_F4(.c1(DAT_WR_E4), .q3(NET00358), .d5(nAD11));
t429 cell_E5(.y3(NET00477), .x5(nDAT_WR));
t406 cell_A5(.c1(NET00442), .r2(NET00444), .q3(NET00443), .r5(GND), .s10(NET00445));
t384 cell_B8(.x1(nDAT_RD), .y3(NET00512), .x5(nDAT_WR));
t389 cell_D35(.x1(WBIT4), .x2(nWCLK), .y3(NET00499), .x4(WBIT2), .y5(NET00497), .x6(NET00499), .x10(NET00500));
t406 cell_I12(.c1(NET00011), .r2(NET00082), .q4(NET00347), .r5(NET00584), .s10(SREG2));
t416 cell_H4(.c1(NET00477), .q3(NET00098), .d5(nAD7));
t416 cell_F5(.c1(DAT_WR_E4), .q3(NET00471), .d5(nAD10));
t417 cell_O7(.x1(NET00139), .y4(NET00147), .x5(NET00140), .x6(NET00596), .x10(OE_RDAT));
t417 cell_J7(.x1(NET00099), .y4(NET00567), .x5(NET00569), .x6(NET00101), .x10(NET00123));
t406 cell_F11(.c1(NET00006), .r2(INIT_073), .q3(SREG5), .q4(nSREG5), .r5(NET00086), .s10(NET00087));
t406 cell_L36(.c1(CRC_CLK1), .r2(CRC_RST3), .q3(CRC15), .q4(nCRC15), .r5(NET00305), .s10(NET00302));
t406 cell_L26(.c1(CRC_CLK1), .r2(CRC_RST0), .q3(NET00066), .q4(NET00068), .r5(NET00065), .s10(NET00067));
t428 cell_K21(.x2(NET00079), .y3(RDINIT1));
t428 cell_K22(.x2(NET00079), .y3(RDINIT0));
t406 cell_O39(.c1(NET00175), .r2(NET00182), .q4(NET00133), .r5(nAD5), .s10(NET00183));
t406 cell_O38(.c1(NET00175), .r2(NET00182), .q4(NET00136), .r5(nAD4), .s10(NET00178));
t406 cell_N34(.c1(CRC_CLK0), .r2(CRC_RST1), .q3(NET00227), .q4(NET00195), .r5(NET00226), .s10(NET00223));
t406 cell_N28(.c1(CRC_CLK0), .r2(CRC_RST2), .q3(NET00234), .q4(NET00193), .r5(NET00587), .s10(NET00588));
t406 cell_L30(.c1(CRC_CLK1), .r2(CRC_RST3), .q3(NET00309), .q4(NET00307), .r5(NET00313), .s10(NET00312));
t406 cell_M30(.c1(CRC_CLK0), .r2(CRC_RST2), .q3(NET00262), .q4(NET00261), .r5(NET00263), .s10(NET00264));
t382 cell_J31(.x1(NET00029), .y2(NET00383), .x3(NET00028), .x4(NET00019), .x5(NET00383), .x6(NET00261), .y8(NET00239));
t406 cell_M26(.c1(CRC_CLK0), .r2(CRC_RST0), .q3(NET00023), .q4(NET00019), .r5(NET00034), .s10(NET00031));
t428 cell_K36(.x2(CRC_RST2), .y3(CRC_RST3));
t406 cell_G12(.c1(NET00011), .r2(NET00082), .q4(NET00050), .r5(NET00047), .s10(SREG4));
t386 cell_C20(.x1(nPLL_A), .y2(PLL_B_DELAYED), .y3(NET00401), .y4(NET00403), .x5(nCLK), .x6(NET00401), .x7(PLL_B0));
t391 cell_B23(.x1(PLL_B0), .x2(nPLL_B), .y3(PLL_B0), .y4(NET00282), .x5(nPLL_C), .x6(PLL_C), .y9(nPLL_6OR7), .x10(PLL_B0));
t406 cell_J12(.c1(STB_P15), .r2(NET00082), .q4(NET00459), .r5(NET00571), .s10(SREG1));
t390 cell_L21(.x1(STB_P09), .y4(NET00077), .x5(MARKER), .x6(nINIT), .y9(NET00079), .x10(nGDR));
t428 cell_K38(.x2(INIT_073), .y3(NET00182));
t406 cell_L35(.c1(nCRC_CLK0), .r2(CRC_RST3), .q3(NET00308), .q4(NET00310), .r5(NET00307), .s10(NET00309));
t406 cell_L29(.c1(nCRC_CLK0), .r2(CRC_RST3), .q3(NET00061), .q4(NET00057), .r5(NET00063), .s10(NET00064));
t428 cell_K39(.x2(NET00219), .y3(NET00175));
t418 cell_J27(.x1(NET00068), .x2(NET00063), .y3(NET00064), .y4(NET00063), .x5(NET00037), .x6(NET00066), .x10(NET00040));
t406 cell_N37(.c1(nCRC_CLK1), .r2(CRC_RST1), .q3(NET00229), .q4(NET00231), .r5(NET00195), .s10(NET00227));
t428 cell_K31(.x2(CRC_CLK0), .y3(CRC_CLK1));
t428 cell_K11(.x2(STB_P15), .y3(CRC_CLK0));
t373 cell_J37(.x1(MODE_R_nW), .x3(nLATCH_TR), .y4(CRC_IN0));
t428 cell_K34(.x2(nCRC_CLK0), .y3(nCRC_CLK1));
t428 cell_E31(.x2(STB_P07), .y3(nCRC_CLK0));
t406 cell_N31(.c1(nCRC_CLK1), .r2(CRC_RST2), .q3(NET00233), .q4(NET00235), .r5(NET00193), .s10(NET00234));
t381 cell_J35(.x1(nCRC15), .y2(CRC_VALID), .x3(NET00301), .x4(NET00385), .x6(NET00307));
t406 cell_N27(.c1(nCRC_CLK1), .r2(CRC_RST0), .q3(NET00591), .q4(NET00590), .r5(NET00240), .s10(NET00607));
t406 cell_G39(.c1(NET00219), .r2(NET00182), .q3(CSR_WM), .r5(nAD9), .s10(NET00380));
t406 cell_M37(.c1(nCRC_CLK1), .r2(CRC_RST1), .q3(NET00258), .q4(NET00256), .r5(NET00254), .s10(NET00253));
t382 cell_O33(.x1(NET00191), .y2(NET00190), .x3(NET00192), .x4(NET00195), .x5(NET00190), .x6(NET00193), .y8(NET00194));
t406 cell_G36(.c1(NET00219), .r2(INIT_F26), .q3(CSR_GDR), .q4(nCSR_GDR), .r5(nAD8), .s10(NET00417));
t370 cell_G34(.y2(NET00417), .x5(nAD8));
t406 cell_M35(.c1(nCRC_CLK1), .r2(CRC_RST1), .q3(NET00260), .q4(NET00259), .r5(NET00261), .s10(NET00262));
t382 cell_N32(.x1(NET00239), .y2(NET00238), .x3(NET00240), .x4(NET00242), .x5(NET00238), .x6(NET00241), .y8(NET00191));
t406 cell_M29(.c1(nCRC_CLK0), .r2(CRC_RST2), .q3(NET00021), .q4(NET00024), .r5(NET00019), .s10(NET00023));
t406 cell_M23(.c1(nCRC_CLK0), .r2(CRC_RST0), .q3(NET00039), .q4(NET00041), .r5(NET00037), .s10(NET00040));
t378 cell_C26(.x1(PLL_H), .y2(NET00407), .x3(nPLL_B), .x5(NET00406));
t406 cell_L37(.c1(nCRC_CLK0), .r2(CRC_RST3), .q3(NET00302), .q4(NET00305), .r5(NET00301), .s10(NET00304));
t406 cell_L27(.c1(nCRC_CLK0), .r2(CRC_RST0), .q3(NET00067), .q4(NET00065), .r5(NET00069), .s10(NET00070));
t406 cell_N35(.c1(nCRC_CLK1), .r2(CRC_RST1), .q3(NET00223), .q4(NET00226), .r5(NET00192), .s10(NET00225));
t382 cell_J30(.x1(NET00194), .y2(NET00384), .x3(NET00068), .x4(NET00069), .x5(NET00384), .x6(NET00062), .y8(NET00385));
t406 cell_N29(.c1(nCRC_CLK1), .r2(CRC_RST2), .q3(NET00588), .q4(NET00587), .r5(NET00241), .s10(NET00589));
t406 cell_L31(.c1(nCRC_CLK0), .r2(CRC_RST3), .q3(NET00312), .q4(NET00313), .r5(NET00062), .s10(NET00059));
t406 cell_M31(.c1(nCRC_CLK1), .r2(CRC_RST2), .q3(NET00264), .q4(NET00263), .r5(NET00028), .s10(NET00026));
t379 cell_H37(.x1(NET00397), .y2(NET00409), .x3(NET00408), .y4(NET00397), .x5(FIN_STB), .x6(NET00409), .x8(NET00410));
t406 cell_N39(.c1(NET00219), .r2(NET00182), .q4(NET00132), .r5(nAD6), .s10(NET00221));
t387 cell_H15(.x1(nBIT_CNT1), .y2(NET00016), .x3(NET00015), .y4(NET00018), .x5(nBIT_CNT2), .x6(NET00017));
t420 cell_J26(.x1(nSREG_Q), .y2(NET00037), .y3(NET00040), .x4(CRC_IN0), .x5(CRC15), .x6(SREG_Q), .x7(NET00037), .x10(nCRC15));
t406 cell_O36(.c1(NET00175), .r2(NET00182), .q4(NET00143), .r5(nAD3), .s10(NET00186));
t378 cell_B26(.x1(NET00405), .y2(NET00415), .x3(NET00407), .x5(PLL_S));
t373 cell_I35(.x1(nLATCH_TR), .x3(nSTB_P03), .y4(NET00387));
t372 cell_J39(.x1(nAD10), .y2(NET00221), .y3(NET00379), .y4(NET00380), .x5(nAD6), .x6(nAD9));
t372 cell_O37(.x1(nAD5), .y2(NET00186), .y3(NET00183), .y4(NET00178), .x5(nAD3), .x6(nAD4));
t406 cell_G35(.c1(RDATA), .r2(INIT_F26), .q4(nGDR), .r5(nCSR_GDR), .s10(CSR_GDR));
t406 cell_O32(.c1(NET00175), .r2(NET00182), .q4(NET00144), .r5(nAD2), .s10(NET00189));
t418 cell_M39(.x1(NET00242), .x2(NET00254), .y3(NET00253), .y4(NET00254), .x5(NET00037), .x6(NET00255), .x10(NET00040));
t406 cell_M27(.c1(nCRC_CLK0), .r2(CRC_RST0), .q3(NET00031), .q4(NET00034), .r5(NET00029), .s10(NET00033));
t378 cell_B24(.x1(NET00407), .y2(NET00406), .x3(PLL_A), .x5(NET00405));
t406 cell_J34(.c1(NET00387), .r2(RDINIT0), .q4(NET00388), .r5(GND), .s10(CRC_VALID));
t379 cell_N23(.x1(NET00592), .y2(NET00595), .x3(NET00593), .y4(NET00592), .x5(INIT_073), .x6(NET00595), .x8(NET00018));

endmodule
//______________________________________________________________________________
//
