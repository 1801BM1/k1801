//
// Copyright (c) 2014-2017 by 1801BM1@gmail.com
//______________________________________________________________________________
//
`timescale 1ns / 100ps

module vp_095
(
   inout[21:0] PIN_nADC,      // CPU Address/Data inverted bus (with gap 18:8)
   inout[7:0]  PIN_nADP,      // PPU Address/Data inverted bus
                              //
   input[2:0]  PIN_RC,        // configuration
   input       PIN_nINITP,    // initialization
   input       PIN_nSYNCC,    //
   input       PIN_nSYNCP,    //
   input       PIN_nA1C_nDLV, // combined with nDLV
   input       PIN_nA1P,      //
   input       PIN_nDLA,      // output address
   input       PIN_nDLD,      // output data
   input       PIN_nCLD,      // output vector
   input       PIN_nWWC,      // CPU writes
   input       PIN_nRDC,      // CPU reads
   input       PIN_nWWP,      // PPU writes
   input       PIN_nRDP,      // PPU reads
   input       PIN_nBSI,      //
                              //
   output      PIN_nCMPC,     //
   output      PIN_nCMPP,     //
   output      PIN_nWD_nRQ,   //
   output      PIN_nBSO       //
);
//______________________________________________________________________________
//
// Autogenerated netlist
//
wire ADP0;
wire ADP1;
wire ADP2;
wire ADP3;
wire ADP4;
wire ADP6;
wire ADP5;
wire ADP7;

wire nADP0;
wire nADP1;
wire nADP2;
wire nADP3;
wire nADP4;
wire nADP5;
wire nADP6;
wire nADP7_0;
wire nADP7;

wire ADC0;
wire ADC1;
wire ADC2;
wire ADC3;
wire ADC4;
wire ADC5;
wire ADC6;
wire ADC7;

wire nADC0;
wire nADC1;
wire nADC2;
wire nADC2_0;
wire nADC3;
wire nADC4;
wire nADC5;
wire nADC6;
wire nADC7;

wire INIT0;
wire INIT1;
wire INIT2;
wire INIT3;
wire INIT4;

wire WC_CSR0;
wire WC_CSR1;
wire WC_DAT;
wire WP_CSR;
wire WP_DAT;
wire nRC_DAT;
wire nRC_CSR;
wire nRP_CSR;
wire nRP_DAT;

wire SA1;
wire SA5;
wire SA6;
wire SA7;

wire nSA0;
wire nSA1;
wire nSA2;
wire nSA3;
wire nSA4;
wire nSA5;

wire RD0;
wire RD1;
wire RD2;
wire RD3;
wire RD4;
wire RD5;
wire RD6;
wire RD7;

wire nRD0;
wire nRD1;
wire nRD2;
wire nRD3;
wire nRD4;
wire nRD5;
wire nRD6;
wire nRD7;

wire nCSR0;
wire nCSR1;
wire nCSR2;
wire nCSR3;
wire nCSR4;
wire nCSR5;
wire nCSR6;
wire nTR_ERR;

wire MRC0;
wire MRC1;
wire MRC3;
wire MRC2;
wire nMRC01;
wire nMRC02;
wire nMRC13;

wire HL0;
wire HL1;
wire HL2;
wire nHL0;
wire nHL1;
wire nHL2;

wire nSYNCC;
wire nSYNCP0;
wire nSYNCP1;
wire nDLD;
wire nDLVL;
wire nDLA0;
wire nDLA1;
wire nDLVH;
wire DLVL;
wire ADCH;
wire nA1P;
wire nA1C;
wire nADC56;
wire nADC47;
wire nCLD;
wire WP_DONE;

wire NET00002, NET00003, NET00004, NET00009, NET00011, NET00014, NET00015, NET00019;
wire NET00020, NET00021, NET00024, NET00026, NET00027, NET00030, NET00031, NET00033;
wire NET00034, NET00035, NET00037, NET00038, NET00039, NET00040, NET00043, NET00044;
wire NET00045, NET00046, NET00047, NET00048, NET00049, NET00051, NET00056, NET00057;
wire NET00058, NET00060, NET00062, NET00064, NET00070, NET00074, NET00075, NET00076;
wire NET00077, NET00078, NET00392, NET00081, NET00083, NET00084, NET00085, NET00087;
wire NET00088, NET00090, NET00092, NET00094, NET00096, NET00097, NET00098, NET00099;
wire NET00100, NET00101, NET00102, NET00104, NET00105, NET00106, NET00108, NET00109;
wire NET00110, NET00112, NET00113, NET00114, NET00115, NET00118, NET00120, NET00121;
wire NET00122, NET00126, NET00127, NET00129, NET00130, NET00131, NET00390, NET00134;
wire NET00135, NET00137, NET00138, NET00141, NET00142, NET00143, NET00144, NET00145;
wire NET00146, NET00147, NET00148, NET00152, NET00153, NET00154, NET00155, NET00156;
wire NET00157, NET00158, NET00159, NET00162, NET00163, NET00166, NET00167, NET00170;
wire NET00172, NET00181, NET00182, NET00183, NET00184, NET00185, NET00186, NET00187;
wire NET00188, NET00189, NET00192, NET00195, NET00196, NET00197, NET00198, NET00199;
wire NET00202, NET00203, NET00204, NET00206, NET00207, NET00208, NET00209, NET00210;
wire NET00212, NET00213, NET00214, NET00215, NET00216, NET00217, NET00218, NET00219;
wire NET00221, NET00222, NET00223, NET00224, NET00225, NET00226, NET00227, NET00228;
wire NET00229, NET00230, NET00231, NET00232, NET00234, NET00235, NET00236, NET00341;
wire NET00239, NET00240, NET00243, NET00244, NET00245, NET00246, NET00247, NET00248;
wire NET00249, NET00250, NET00251, NET00253, NET00254, NET00255, NET00256, NET00257;
wire NET00258, NET00259, NET00260, NET00261, NET00262, NET00263, NET00264, NET00265;
wire NET00266, NET00267, NET00268, NET00269, NET00270, NET00271, NET00272, NET00273;
wire NET00274, NET00275, NET00276, NET00278, NET00279, NET00281, NET00282, NET00283;
wire NET00284, NET00285, NET00286, NET00287, NET00290, NET00295, NET00297, NET00299;
wire NET00300, NET00298, NET00302, NET00303, NET00301, NET00304, NET00305, NET00307;
wire NET00308, NET00309, NET00310, NET00311, NET00312, NET00314, NET00315, NET00316;
wire NET00319, NET00320, NET00321, NET00323, NET00324, NET00322, NET00391, NET00328;
wire NET00329, NET00331, NET00332, NET00330, NET00333, NET00334, NET00335, NET00338;
wire NET00339, NET00340, NET00342, NET00355, NET00343, NET00344, NET00345, NET00347;
wire NET00348, NET00346, NET00349, NET00350, NET00351, NET00353, NET00354, NET00358;
wire NET00356, NET00357, NET00359, NET00361, NET00360, NET00362, NET00377, NET00364;
wire NET00365, NET00363, NET00366, NET00367, NET00368, NET00370, NET00371, NET00372;
wire NET00373, NET00374, NET00376, NET00385, NET00375, NET00379, NET00381, NET00382;
wire NET00383, NET00384, NET00387, NET00388;

//______________________________________________________________________________
//
// Autogenerated cell instantiations
//
assign PIN_nADC[18:8] = 11'bzzzzzzzzzzz;

tOUTPUT cell_PIN20(.x1(NET00162), .y1(PIN_nCMPC));
tOUTPUT cell_PIN22(.x1(NET00254), .y1(PIN_nCMPP));
tOUTPUT cell_PIN23(.x1(NET00253), .y1(PIN_nWD_nRQ));
tOUTPUT cell_PIN25(.x1(NET00245), .y1(PIN_nBSO));

tOUTPUT_OC cell_PIN6_OC (.x1(NET00060), .y1(PIN_nADC[0]));
tOUTPUT_OC cell_PIN7_OC (.x1(NET00330), .y1(PIN_nADC[1]));
tOUTPUT_OC cell_PIN8_OC (.x1(NET00248), .y1(PIN_nADC[2]));
tOUTPUT_OC cell_PIN9_OC (.x1(NET00363), .y1(PIN_nADC[3]));
tOUTPUT_OC cell_PIN10_OC(.x1(NET00246), .y1(PIN_nADC[4]));
tOUTPUT_OC cell_PIN11_OC(.x1(NET00240), .y1(PIN_nADC[5]));
tOUTPUT_OC cell_PIN12_OC(.x1(NET00083), .y1(PIN_nADC[6]));
tOUTPUT_OC cell_PIN13_OC(.x1(NET00223), .y1(PIN_nADC[7]));
tOUTPUT_OC cell_PIN17_OC(.x1(NET00046), .y1(PIN_nADC[19]));
tOUTPUT_OC cell_PIN18_OC(.x1(NET00048), .y1(PIN_nADC[20]));
tOUTPUT_OC cell_PIN19_OC(.x1(NET00045), .y1(PIN_nADC[21]));

tOUTPUT_OC cell_PIN35_OC(.x1(NET00085), .y1(PIN_nADP[0]));
tOUTPUT_OC cell_PIN34_OC(.x1(NET00154), .y1(PIN_nADP[1]));
tOUTPUT_OC cell_PIN33_OC(.x1(NET00182), .y1(PIN_nADP[2]));
tOUTPUT_OC cell_PIN32_OC(.x1(NET00262), .y1(PIN_nADP[3]));
tOUTPUT_OC cell_PIN31_OC(.x1(NET00274), .y1(PIN_nADP[4]));
tOUTPUT_OC cell_PIN30_OC(.x1(NET00251), .y1(PIN_nADP[5]));
tOUTPUT_OC cell_PIN29_OC(.x1(NET00346), .y1(PIN_nADP[6]));
tOUTPUT_OC cell_PIN28_OC(.x1(NET00298), .y1(PIN_nADP[7]));

tINPUT cell_PIN6 (.y2(NET00094), .x1(PIN_nADC[0]));
tINPUT cell_PIN7 (.y2(NET00090), .x1(PIN_nADC[1]));
tINPUT cell_PIN8 (.y2(NET00088), .x1(PIN_nADC[2]));
tINPUT cell_PIN9 (.y2(NET00101), .x1(PIN_nADC[3]));
tINPUT cell_PIN10(.y2(NET00392), .x1(PIN_nADC[4]));
tINPUT cell_PIN11(.y2(NET00316), .x1(PIN_nADC[5]));
tINPUT cell_PIN12(.y2(NET00314), .x1(PIN_nADC[6]));
tINPUT cell_PIN13(.y2(NET00315), .x1(PIN_nADC[7]));
tINPUT cell_PIN17(.y1(NET00228), .x1(PIN_nADC[19]));
tINPUT cell_PIN18(.y1(NET00230), .x1(PIN_nADC[20]));
tINPUT cell_PIN19(.y1(NET00229), .x1(PIN_nADC[21]));

tINPUT cell_PIN35(.y2(NET00092), .x1(PIN_nADP[0]));
tINPUT cell_PIN34(.y2(NET00087), .x1(PIN_nADP[1]));
tINPUT cell_PIN33(.y2(NET00105), .x1(PIN_nADP[2]));
tINPUT cell_PIN32(.y2(NET00102), .x1(PIN_nADP[3]));
tINPUT cell_PIN31(.y2(NET00100), .x1(PIN_nADP[4]));
tINPUT cell_PIN30(.y2(NET00099), .x1(PIN_nADP[5]));
tINPUT cell_PIN29(.y2(NET00260), .x1(PIN_nADP[6]));
tINPUT cell_PIN28(.y2(NET00261), .x1(PIN_nADP[7]));

tINPUT cell_PIN2 (.y2(NET00051), .x1(PIN_RC[0]));
tINPUT cell_PIN1 (.y1(NET00113), .x1(PIN_RC[1]));
tINPUT cell_PIN41(.y1(NET00114), .x1(PIN_RC[2]));

tINPUT cell_PIN37(.y2(NET00098), .x1(PIN_nINITP));
tINPUT cell_PIN38(.y1(NET00035), .x1(PIN_nSYNCP));
tINPUT cell_PIN4 (.y1(nSYNCC),   .x1(PIN_nSYNCC));

tINPUT cell_PIN5 (.y1(NET00097), .x1(PIN_nDLA));
tINPUT cell_PIN14(.y1(NET00081), .x1(PIN_nDLD));
tINPUT cell_PIN36(.y1(NET00096), .x1(PIN_nCLD));
tINPUT cell_PIN15(.y1(NET00322), .x1(PIN_nWWC));
tINPUT cell_PIN16(.y1(NET00301), .x1(PIN_nRDC));
tINPUT cell_PIN27(.y1(NET00217), .x1(PIN_nWWP));
tINPUT cell_PIN26(.y1(NET00390), .x1(PIN_nRDP));

tINPUT cell_PIN40(.y2(NET00375), .x1(PIN_nA1P));
tINPUT cell_PIN3 (.y2(NET00122), .x1(PIN_nA1C_nDLV));
tINPUT cell_PIN39(.y2(NET00106), .x1(PIN_nBSI));

t408 cell_A22(.q2(RD7), .q3(nRD7), .r5(NET00192), .s10(NET00195));
t390 cell_O35(.x1(RD0), .y4(NET00126), .x5(HL1), .x6(SA5), .y9(NET00127), .x10(HL1));
t376 cell_A21(.x1(nRP_DAT), .x3(nRD7), .y4(NET00297), .x6(nRC_DAT), .x8(nRD7), .y9(NET00224));
t428 cell_E39(.x2(NET00261), .y3(ADP7));
t408 cell_C22(.q2(RD6), .q3(nRD6), .r5(NET00167), .s10(NET00166));
t428 cell_E2(.x2(NET00316), .y3(ADC5));
t390 cell_C35(.x1(RD7), .y4(NET00343), .x5(nHL2), .x6(RD6), .y9(NET00344), .x10(nHL2));
t373 cell_C28(.x1(nCSR6), .x3(nRP_CSR), .y4(NET00283));
t428 cell_K12(.x2(INIT1), .y3(INIT4));
t373 cell_N0(.x1(NET00375), .x3(nHL0), .y4(NET00312));
t387 cell_O0(.x1(nHL0), .y2(nDLVL), .x3(nHL0), .y4(nDLVH), .x5(NET00122), .x6(NET00122));
t373 cell_M28(.x1(nCSR2), .x3(nRP_CSR), .y4(NET00002));
t379 cell_N14(.x1(nSA1), .y2(SA1), .x3(NET00351), .y4(nSA1), .x5(INIT2), .x6(SA1), .x8(NET00353));
t376 cell_N21(.x1(nRP_DAT), .x3(nRD1), .y4(NET00153), .x6(nRC_DAT), .x8(nRD1), .y9(NET00331));
t378 cell_I33(.x1(NET00273), .y2(NET00274), .x3(NET00137), .x5(NET00142));
t377 cell_J37(.x1(NET00267), .y2(NET00267), .x3(nMRC13), .y4(NET00268), .x5(ADP2), .x6(nMRC02), .x8(ADP2), .y9(NET00269));
t391 cell_J38(.x1(ADP6), .x2(ADP1), .y3(NET00256), .y4(NET00257), .x5(NET00255), .x6(ADP2), .y9(NET00258), .x10(ADP3));
t378 cell_J33(.x1(NET00183), .y2(NET00262), .x3(NET00104), .x5(NET00108));
t408 cell_A24(.q3(nTR_ERR), .r5(NET00188), .s10(NET00299));
t379 cell_B4(.x1(NET00365), .y2(nA1C), .x3(NET00308), .y4(NET00365), .x5(INIT0), .x6(nA1C), .x8(NET00310));
t408 cell_C26(.q3(nCSR6), .r5(NET00281), .s10(NET00282));
t428 cell_E4(.x2(NET00392), .y3(ADC4));
t380 cell_D0(.x1(NET00076), .y2(NET00227), .y3(NET00226), .x4(NET00227), .x5(MRC3), .x6(nADC2_0));
t371 cell_C37(.x1(ADP7), .y3(nADP7), .y4(nADP6), .x6(ADP6));
t380 cell_J2(.x1(nADC2_0), .y2(NET00368), .y3(NET00321), .x4(NET00368), .x5(MRC1), .x6(ADC3));
t389 cell_H2(.x1(NET00235), .x2(ADP7), .y3(NET00020), .x4(nMRC02), .y5(NET00234), .x6(ADCH), .x10(NET00236));
t376 cell_I16(.x1(nADP5), .x3(nDLD), .y4(NET00239), .x6(nADP4), .x8(nDLD), .y9(NET00324));
t381 cell_I6(.x1(NET00323), .y2(NET00246), .x3(NET00324), .x4(NET00319), .x6(NET00143));
t408 cell_I26(.q3(nCSR4), .r5(NET00144), .s10(NET00145));
t379 cell_O12(.x1(NET00341), .y2(NET00340), .x3(nSYNCP1), .y4(NET00341), .x5(NET00338), .x6(NET00340), .x8(ADP0));
t373 cell_I28(.x1(nCSR4), .x3(nRP_CSR), .y4(NET00137));
t428 cell_K35(.x2(NET00092), .y3(ADP0));
t378 cell_M33(.x1(NET00181), .y2(NET00182), .x3(NET00002), .x5(NET00014));
t378 cell_N33(.x1(NET00152), .y2(NET00154), .x3(NET00155), .x5(NET00153));
t379 cell_C10(.x1(NET00156), .y2(NET00159), .x3(INIT1), .y4(NET00156), .x5(NET00157), .x6(NET00159), .x8(nSYNCP0));
t383 cell_H6(.x1(DLVL), .y2(NET00240), .x3(NET00239), .x4(NET00221), .x5(NET00064), .x6(NET00203));
t428 cell_E12(.x2(WP_DAT), .y3(NET00031));
t371 cell_D4(.x1(ADC7), .y3(nADC7), .y4(nADC6), .x6(ADC6));
t381 cell_D6(.x1(NET00057), .y2(NET00223), .x3(NET00134), .x4(NET00225), .x6(NET00224));
t428 cell_E6(.x2(WC_DAT), .y3(NET00033));
t379 cell_J10(.x1(NET00372), .y2(NET00376), .x3(INIT2), .y4(NET00372), .x5(NET00373), .x6(NET00376), .x8(nSYNCP1));
t379 cell_M10(.x1(NET00357), .y2(NET00362), .x3(INIT2), .y4(NET00357), .x5(NET00361), .x6(NET00362), .x8(nSYNCP1));
t408 cell_J26(.q3(nCSR3), .r5(NET00120), .s10(NET00121));
t379 cell_O14(.x1(nSA0), .y2(NET00339), .x3(NET00338), .y4(nSA0), .x5(INIT2), .x6(NET00339), .x8(NET00340));
t428 cell_K37(.x2(NET00087), .y3(ADP1));
t428 cell_K38(.x2(NET00105), .y3(ADP2));
t379 cell_B12(.x1(NET00185), .y2(NET00186), .x3(nSYNCP0), .y4(NET00185), .x5(NET00184), .x6(NET00186), .x8(ADP7));
t377 cell_G9(.x1(HL0), .y2(NET00056), .x3(NET00078), .y4(WP_DONE), .x5(NET00077), .x6(HL0), .x8(nRC_CSR), .y9(NET00077));
t376 cell_G6(.x1(nDLA1), .x3(NET00062), .y4(NET00044), .x6(nSA5), .x8(nDLA0), .y9(NET00064));
t418 cell_D26(.x1(nHL2), .x2(NET00021), .y3(NET00271), .y4(NET00253), .x5(NET00270), .x6(HL1), .x10(NET00271));
t428 cell_E25(.x2(nHL0), .y3(nHL1));
t376 cell_D16(.x1(nADP7), .x3(nDLD), .y4(NET00134), .x6(nADP6), .x8(nDLD), .y9(NET00135));
t428 cell_E16(.x2(INIT0), .y3(INIT3));
t379 cell_N10(.x1(NET00351), .y2(NET00355), .x3(INIT2), .y4(NET00351), .x5(NET00354), .x6(NET00355), .x8(nSYNCP1));
t379 cell_O10(.x1(NET00338), .y2(NET00342), .x3(INIT2), .y4(NET00338), .x5(NET00341), .x6(NET00342), .x8(nSYNCP1));
t373 cell_J28(.x1(nCSR3), .x3(nRP_CSR), .y4(NET00104));
t428 cell_K24(.x2(NET00049), .y3(WC_CSR1));
t379 cell_J14(.x1(nSA3), .y2(NET00377), .x3(NET00372), .y4(nSA3), .x5(INIT2), .x6(NET00377), .x8(NET00374));
t380 cell_L4(.x1(ADC3), .y2(NET00244), .y3(NET00243), .x4(NET00244), .x5(MRC0), .x6(ADC2));
t389 cell_C2(.x1(NET00037), .x2(NET00039), .y3(NET00038), .x4(nADC56), .y5(NET00037), .x6(ADCH), .x10(NET00040));
t390 cell_M35(.x1(RD2), .y4(NET00146), .x5(HL1), .x6(RD1), .y9(NET00148), .x10(HL1));
t428 cell_K31(.x2(NET00098), .y3(INIT0));
t379 cell_B14(.x1(NET00189), .y2(SA7), .x3(NET00184), .y4(NET00189), .x5(INIT1), .x6(SA7), .x8(NET00186));
t379 cell_C12(.x1(NET00157), .y2(NET00158), .x3(nSYNCP0), .y4(NET00157), .x5(NET00156), .x6(NET00158), .x8(ADP6));
t379 cell_G12(.x1(NET00027), .y2(NET00026), .x3(nSYNCP0), .y4(NET00027), .x5(NET00024), .x6(NET00026), .x8(ADP5));
t379 cell_G10(.x1(NET00024), .y2(NET00030), .x3(INIT1), .y4(NET00024), .x5(NET00027), .x6(NET00030), .x8(nSYNCP0));
t428 cell_E38(.x2(NET00260), .y3(ADP6));
t428 cell_E32(.x2(HL0), .y3(HL1));
t387 cell_D28(.x1(WP_DONE), .y2(NET00272), .x3(NET00272), .y4(NET00270), .x5(ADP5), .x6(nCSR6));
t376 cell_D30(.x1(nADC7), .x3(nCLD), .y4(NET00347), .x6(nADC6), .x8(nCLD), .y9(NET00345));
t379 cell_M14(.x1(nSA2), .y2(NET00358), .x3(NET00357), .y4(nSA2), .x5(INIT2), .x6(NET00358), .x8(NET00359));
t429 cell_K26(.y3(HL0), .x5(NET00051));
t376 cell_L2(.x1(MRC1), .x3(MRC0), .y4(nMRC01), .x6(MRC0), .x8(MRC2), .y9(nMRC02));
t428 cell_K33(.x2(NET00096), .y3(nCLD));
t372 cell_M37(.x1(ADP2), .y2(nADP0), .y3(nADP2), .y4(nADP1), .x5(ADP0), .x6(ADP1));
t419 cell_B16(.x1(WP_CSR), .y2(NET00188), .x4(INIT0), .x5(nADP7), .x6(nHL0), .x10(NET00033));
t379 cell_G14(.x1(nSA5), .y2(SA5), .x3(NET00024), .y4(nSA5), .x5(INIT1), .x6(SA5), .x8(NET00026));
t379 cell_I10(.x1(NET00382), .y2(NET00383), .x3(INIT1), .y4(NET00382), .x5(NET00381), .x6(NET00383), .x8(nSYNCP0));
t381 cell_D35(.x1(NET00343), .y2(NET00300), .x3(NET00344), .x4(nDLA1), .x6(NET00290));
t428 cell_E35(.x2(NET00100), .y3(ADP4));
t428 cell_E37(.x2(NET00099), .y3(ADP5));
t408 cell_I22(.q2(RD4), .q3(nRD4), .r5(NET00138), .s10(NET00141));
t376 cell_I21(.x1(nRP_DAT), .x3(nRD4), .y4(NET00142), .x6(nRC_DAT), .x8(nRD4), .y9(NET00143));
t428 cell_K28(.x2(NET00035), .y3(nSYNCP1));
t417 cell_J18(.x1(NET00332), .y4(NET00112), .x5(ADP3), .x6(NET00333), .x10(ADC3));
t390 cell_I35(.x1(RD4), .y4(NET00265), .x5(HL1), .x6(RD3), .y9(NET00266), .x10(HL1));
t376 cell_N30(.x1(nADC1), .x3(nCLD), .y4(NET00152), .x6(nADC0), .x8(nCLD), .y9(NET00130));
t417 cell_B18(.x1(NET00031), .y4(NET00195), .x5(ADP7), .x6(NET00033), .x10(ADC7));
t379 cell_I12(.x1(NET00381), .y2(NET00384), .x3(nSYNCP0), .y4(NET00381), .x5(NET00382), .x6(NET00384), .x8(ADP4));
t429 cell_E7(.y3(nRC_CSR), .x5(NET00305));
t428 cell_E1(.x2(NET00314), .y3(ADC6));
t390 cell_F2(.x1(ADC5), .y4(nADC56), .x5(ADC6), .x6(ADC4), .y9(nADC47), .x10(ADC7));
t429 cell_E28(.y3(nRP_CSR), .x5(NET00259));
t376 cell_J21(.x1(nRP_DAT), .x3(nRD3), .y4(NET00108), .x6(nRC_DAT), .x8(nRD3), .y9(NET00109));
t379 cell_N12(.x1(NET00354), .y2(NET00353), .x3(nSYNCP1), .y4(NET00354), .x5(NET00351), .x6(NET00353), .x8(ADP1));
t428 cell_K16(.x2(WP_DAT), .y3(NET00332));
t408 cell_M26(.q3(nCSR2), .r5(NET00003), .s10(NET00004));
t419 cell_J19(.x1(NET00332), .y2(NET00110), .x4(INIT4), .x5(nADP3), .x6(NET00333), .x10(nADC3));
t381 cell_J35(.x1(NET00263), .y2(NET00264), .x3(NET00265), .x4(nDLA1), .x6(NET00266));
t376 cell_I37(.x1(NET00275), .x3(NET00257), .y4(NET00276), .x6(NET00268), .x8(NET00269), .y9(NET00275));
t408 cell_H28(.q3(nCSR5), .r5(NET00170), .s10(NET00172));
t379 cell_I14(.x1(nSA4), .y2(NET00385), .x3(NET00382), .y4(nSA4), .x5(INIT1), .x6(NET00385), .x8(NET00384));
t408 cell_G22(.q2(RD5), .q3(nRD5), .r5(NET00204), .s10(NET00034));
t392 cell_F35(.x1(NET00264), .x3(NET00300), .y4(NET00245), .x5(NET00147));
t428 cell_K1(.x2(NET00090), .y3(ADC1));
t381 cell_F37(.x1(ADP3), .y2(NET00255), .x3(ADP4), .x4(ADP7), .x6(ADP5));
t428 cell_K0(.x2(NET00094), .y3(ADC0));
t376 cell_F8(.x1(nDLA1), .x3(NET00356), .y4(NET00225), .x6(nDLA1), .x8(NET00295), .y9(NET00367));
t429 cell_E33(.y3(nHL2), .x5(HL0));
t390 cell_F38(.x1(ADP5), .y4(NET00286), .x5(ADP4), .x6(ADP7), .y9(NET00284), .x10(ADP6));
t383 cell_F6(.x1(DLVL), .y2(NET00083), .x3(NET00135), .x4(NET00058), .x5(NET00367), .x6(NET00279));
t419 cell_M19(.x1(NET00332), .y2(NET00009), .x4(INIT4), .x5(nADP2), .x6(NET00333), .x10(nADC2));
t376 cell_M16(.x1(nADP3), .x3(nDLD), .y4(NET00360), .x6(nADP2), .x8(nDLD), .y9(NET00249));
t417 cell_O18(.x1(NET00332), .y4(NET00334), .x5(ADP0), .x6(NET00333), .x10(ADC0));
t382 cell_I2(.x1(NET00243), .y2(NET00039), .x3(NET00074), .x4(NET00321), .x5(ADP6), .x6(NET00226), .y8(NET00235));
t417 cell_G18(.x1(NET00031), .y4(NET00034), .x5(ADP5), .x6(NET00033), .x10(ADC5));
t383 cell_H38(.x1(ADP0), .y2(NET00285), .x3(NET00258), .x4(NET00256), .x5(NET00284), .x6(NET00286));
t379 cell_J4(.x1(ADC0), .y2(NET00236), .x3(ADC1), .y4(nMRC13), .x5(ADC3), .x6(MRC1), .x8(MRC3));
t417 cell_G28(.x1(NET00198), .y4(NET00172), .x5(ADC5), .x6(WP_DONE), .x10(ADP5));
t428 cell_K2(.x2(NET00088), .y3(ADC2));
t419 cell_C20(.x1(NET00031), .y2(NET00204), .x4(INIT4), .x5(nADP5), .x6(NET00033), .x10(nADC5));
t376 cell_M8(.x1(nDLA0), .x3(nSA2), .y4(NET00250), .x6(nSA1), .x8(nDLA0), .y9(NET00328));
t408 cell_O26(.q3(nCSR0), .r5(NET00379), .s10(NET00197));
t373 cell_O28(.x1(nCSR0), .x3(nRP_CSR), .y4(NET00131));
t429 cell_E8(.y3(nRC_DAT), .x5(NET00304));
t376 cell_A0(.x1(NET00301), .x3(NET00302), .y4(NET00304), .x6(NET00301), .x8(NET00303), .y9(NET00305));
t419 cell_B19(.x1(NET00031), .y2(NET00192), .x4(INIT4), .x5(nADP7), .x6(NET00033), .x10(nADC7));
t376 cell_B0(.x1(NET00322), .x3(NET00302), .y4(WC_DAT), .x6(NET00322), .x8(NET00303), .y9(NET00049));
t429 cell_E10(.y3(NET00078), .x5(WP_CSR));
t376 cell_C21(.x1(nRP_DAT), .x3(nRD6), .y4(NET00278), .x6(nRC_DAT), .x8(nRD6), .y9(NET00279));
t419 cell_C19(.x1(NET00031), .y2(NET00167), .x4(INIT4), .x5(nADP6), .x6(NET00033), .x10(nADC6));
t377 cell_I4(.x1(nMRC13), .y2(DLVL), .x3(nDLVL), .y4(NET00247), .x5(nDLVL), .x6(nDLVL), .x8(nMRC01), .y9(NET00323));
t376 cell_A18(.x1(NET00390), .x3(NET00218), .y4(NET00084), .x6(NET00390), .x8(NET00219), .y9(NET00259));
t398 cell_I24(.x1(WC_CSR0), .y2(NET00144), .x4(INIT3), .x5(nADC4), .x6(ADC4), .y9(NET00145), .x10(WC_CSR0));
t376 cell_M21(.x1(nRP_DAT), .x3(nRD2), .y4(NET00014), .x6(nRC_DAT), .x8(nRD2), .y9(NET00015));
t375 cell_A2(.x1(NET00215), .y2(NET00303), .y3(NET00302), .x4(nA1C), .x5(NET00303), .x6(ADC2), .y9(nADC2_0));
t429 cell_E26(.y3(HL2), .x5(nHL0));
t379 cell_A4(.x1(NET00308), .y2(NET00309), .x3(INIT0), .y4(NET00308), .x5(NET00307), .x6(NET00309), .x8(nSYNCC));
t417 cell_B24(.x1(RD7), .y4(NET00062), .x5(nHL1), .x6(RD4), .x10(HL2));
t429 cell_E14(.y3(nRP_DAT), .x5(NET00084));
t398 cell_C24(.x1(WC_CSR1), .y2(NET00281), .x4(INIT3), .x5(nADC6), .x6(ADC6), .y9(NET00282), .x10(WC_CSR1));
t417 cell_C18(.x1(NET00031), .y4(NET00166), .x5(ADP6), .x6(NET00033), .x10(ADC6));
t376 cell_N16(.x1(nADP1), .x3(nDLD), .y4(NET00329), .x6(nADP0), .x8(nDLD), .y9(NET00350));
t417 cell_B26(.x1(RD6), .y4(NET00231), .x5(nHL1), .x6(RD3), .x10(HL2));
t376 cell_D8(.x1(nDLA1), .x3(NET00231), .y4(NET00047), .x6(nDLA1), .x8(NET00232), .y9(NET00043));
t376 cell_I8(.x1(nDLA0), .x3(nSA4), .y4(NET00319), .x6(nSA3), .x8(nDLA0), .y9(NET00320));
t379 cell_A6(.x1(NET00307), .y2(NET00310), .x3(nSYNCC), .y4(NET00307), .x5(NET00308), .x6(NET00310), .x8(nDLVH));
t398 cell_J24(.x1(WC_CSR1), .y2(NET00120), .x4(INIT3), .x5(nADC3), .x6(ADC3), .y9(NET00121), .x10(WC_CSR1));
t379 cell_A8(.x1(NET00206), .y2(NET00311), .x3(nSYNCP0), .y4(NET00206), .x5(NET00207), .x6(NET00311), .x8(NET00312));
t372 cell_M2(.x1(ADC2), .y2(nADC0), .y3(nADC2), .y4(nADC1), .x5(ADC0), .x6(ADC1));
t376 cell_A16(.x1(NET00217), .x3(NET00218), .y4(WP_DAT), .x6(NET00217), .x8(NET00219), .y9(WP_CSR));
t384 cell_B33(.x1(ADP7), .y3(NET00299), .x5(WP_CSR));
t417 cell_B28(.x1(RD5), .y4(NET00232), .x5(nHL1), .x6(RD2), .x10(HL2));
t377 cell_O2(.x1(NET00113), .y2(NET00118), .x3(NET00118), .y4(MRC2), .x5(NET00114), .x6(NET00118), .x8(NET00115), .y9(MRC3));
t378 cell_M6(.x1(NET00329), .y2(NET00330), .x3(NET00331), .x5(NET00328));
t376 cell_C8(.x1(nTR_ERR), .x3(nRC_CSR), .y4(NET00057), .x6(nCSR6), .x8(NET00056), .y9(NET00058));
t379 cell_C14(.x1(NET00163), .y2(SA6), .x3(NET00156), .y4(NET00163), .x5(INIT1), .x6(SA6), .x8(NET00158));
t379 cell_A14(.x1(NET00209), .y2(NET00216), .x3(INIT0), .y4(NET00209), .x5(NET00210), .x6(NET00216), .x8(nSYNCC));
t379 cell_A13(.x1(NET00214), .y2(NET00215), .x3(NET00209), .y4(NET00214), .x5(INIT0), .x6(NET00215), .x8(NET00212));
t417 cell_C30(.x1(SA7), .y4(NET00356), .x5(nHL1), .x6(RD1), .x10(HL2));
t380 cell_G0(.x1(ADC2), .y2(NET00075), .y3(NET00074), .x4(NET00075), .x5(MRC2), .x6(NET00076));
t390 cell_G35(.x1(RD5), .y4(NET00290), .x5(nHL2), .x6(NET00106), .y9(NET00263), .x10(HL1));
t378 cell_C33(.x1(NET00287), .y2(NET00251), .x3(NET00222), .x5(NET00202));
t398 cell_N24(.x1(WC_CSR0), .y2(NET00387), .x4(INIT3), .x5(nADC1), .x6(ADC1), .y9(NET00388), .x10(WC_CSR0));
t408 cell_J22(.q2(RD3), .q3(nRD3), .r5(NET00110), .s10(NET00112));
t372 cell_G37(.x1(ADP5), .y2(nADP3), .y3(nADP5), .y4(nADP4), .x5(ADP3), .x6(ADP4));
t408 cell_N22(.q2(RD1), .q3(nRD1), .r5(NET00348), .s10(NET00349));
t379 cell_B8(.x1(NET00366), .y2(nA1P), .x3(NET00207), .y4(NET00366), .x5(INIT0), .x6(nA1P), .x8(NET00311));
t379 cell_B10(.x1(NET00184), .y2(NET00187), .x3(INIT1), .y4(NET00184), .x5(NET00185), .x6(NET00187), .x8(nSYNCP0));
t428 cell_K39(.x2(NET00102), .y3(ADP3));
t372 cell_G4(.x1(ADC5), .y2(nADC3), .y3(nADC5), .y4(nADC4), .x5(ADC3), .x6(ADC4));
t379 cell_D2(.x1(NET00229), .y2(ADCH), .x3(NET00230), .y4(NET00040), .x5(NET00228), .x6(ADC4), .x8(ADC7));
t376 cell_F28(.x1(NET00056), .x3(nCSR5), .y4(NET00221), .x6(nCSR5), .x8(nRP_CSR), .y9(NET00222));
t379 cell_M12(.x1(NET00361), .y2(NET00359), .x3(nSYNCP1), .y4(NET00361), .x5(NET00357), .x6(NET00359), .x8(ADP2));
t381 cell_J6(.x1(DLVL), .y2(NET00363), .x3(NET00360), .x4(NET00320), .x6(NET00109));
t428 cell_K25(.x2(NET00049), .y3(WC_CSR0));
t376 cell_G21(.x1(nRP_DAT), .x3(nRD5), .y4(NET00202), .x6(nRC_DAT), .x8(nRD5), .y9(NET00203));
t373 cell_N28(.x1(nCSR1), .x3(nRP_CSR), .y4(NET00155));
t381 cell_L6(.x1(NET00247), .y2(NET00248), .x3(NET00249), .x4(NET00250), .x6(NET00015));
t383 cell_N35(.x1(NET00146), .y2(NET00147), .x3(NET00126), .x4(NET00148), .x5(nDLA1), .x6(NET00127));
t428 cell_K32(.x2(NET00098), .y3(INIT1));
t428 cell_K30(.x2(NET00035), .y3(nSYNCP0));
t378 cell_O33(.x1(NET00130), .y2(NET00085), .x3(NET00131), .x5(NET00129));
t417 cell_H37(.x1(HL0), .y4(NET00254), .x5(NET00285), .x6(nHL2), .x10(NET00276));
t376 cell_H30(.x1(nADC5), .x3(nCLD), .y4(NET00287), .x6(nADC4), .x8(nCLD), .y9(NET00273));
t376 cell_M30(.x1(nADC3), .x3(nCLD), .y4(NET00183), .x6(nADC2), .x8(nCLD), .y9(NET00181));
t379 cell_B30(.x1(NET00347), .y2(NET00298), .x3(NET00364), .y4(NET00364), .x5(NET00297), .x6(nTR_ERR), .x8(nRP_CSR));
t417 cell_G30(.x1(SA6), .y4(NET00295), .x5(nHL1), .x6(RD0), .x10(HL2));
t372 cell_C6(.x1(NET00044), .y2(NET00046), .y3(NET00045), .y4(NET00048), .x5(NET00043), .x6(NET00047));
t381 cell_G2(.x1(NET00234), .y2(NET00070), .x3(nADC2_0), .x4(nADC47), .x6(nADC56));
t378 cell_D33(.x1(NET00345), .y2(NET00346), .x3(NET00283), .x5(NET00278));
t375 cell_H8(.x1(NET00391), .y2(NET00219), .y3(NET00218), .x4(nA1P), .x5(NET00219), .x6(ADC3), .y9(NET00076));
t428 cell_E0(.x2(NET00315), .y3(ADC7));
t379 cell_J12(.x1(NET00373), .y2(NET00374), .x3(nSYNCP1), .y4(NET00373), .x5(NET00372), .x6(NET00374), .x8(ADP3));
t428 cell_K15(.x2(WC_DAT), .y3(NET00333));
t417 cell_M18(.x1(NET00332), .y4(NET00011), .x5(ADP2), .x6(NET00333), .x10(ADC2));
t417 cell_N18(.x1(NET00332), .y4(NET00349), .x5(ADP1), .x6(NET00333), .x10(ADC1));
t373 cell_J16(.x1(HL0), .x3(ADC1), .y4(NET00213));
t408 cell_N26(.q3(nCSR1), .r5(NET00387), .s10(NET00388));
t417 cell_I18(.x1(NET00031), .y4(NET00141), .x5(ADP4), .x6(NET00033), .x10(ADC4));
t419 cell_I19(.x1(NET00031), .y2(NET00138), .x4(INIT4), .x5(nADP4), .x6(NET00033), .x10(nADC4));
t428 cell_K27(.x2(NET00051), .y3(nHL0));
t419 cell_N19(.x1(NET00332), .y2(NET00348), .x4(INIT4), .x5(nADP1), .x6(NET00333), .x10(nADC1));
t419 cell_O19(.x1(NET00332), .y2(NET00335), .x4(INIT4), .x5(nADP0), .x6(NET00333), .x10(nADC0));
t377 cell_G24(.x1(NET00196), .y2(NET00196), .x3(nHL0), .y4(NET00198), .x5(WC_CSR1), .x6(HL0), .x8(NET00197), .y9(NET00199));
t421 cell_G26(.x1(WP_DONE), .y2(NET00170), .x3(NET00199), .x4(INIT3), .x5(nADP5), .x6(NET00198), .x10(nADC5));
t428 cell_K8(.x2(NET00081), .y3(nDLD));
t428 cell_K10(.x2(INIT0), .y3(INIT2));
t428 cell_K4(.x2(NET00101), .y3(ADC3));
t428 cell_K7(.x2(NET00097), .y3(nDLA1));
t428 cell_K6(.x2(NET00097), .y3(nDLA0));
t408 cell_O22(.q2(RD0), .q3(nRD0), .r5(NET00335), .s10(NET00334));
t379 cell_A10(.x1(NET00207), .y2(NET00208), .x3(INIT0), .y4(NET00207), .x5(NET00206), .x6(NET00208), .x8(nSYNCP0));
t379 cell_A12(.x1(NET00210), .y2(NET00212), .x3(nSYNCC), .y4(NET00210), .x5(NET00209), .x6(NET00212), .x8(NET00213));
t377 cell_O4(.x1(NET00113), .y2(NET00115), .x3(NET00114), .y4(MRC0), .x5(NET00113), .x6(NET00115), .x8(NET00114), .y9(MRC1));
t379 cell_G16(.x1(ADP6), .y2(NET00019), .x3(nMRC13), .y4(NET00021), .x5(nADP7_0), .x6(NET00019), .x8(NET00020));
t378 cell_N6(.x1(NET00350), .y2(NET00060), .x3(NET00371), .x5(NET00370));
t418 cell_C16(.x1(NET00070), .x2(ADP7), .y3(nADP7_0), .y4(NET00162), .x5(HL1), .x6(nHL2), .x10(NET00038));
t398 cell_M24(.x1(WC_CSR0), .y2(NET00003), .x4(INIT3), .x5(nADC2), .x6(ADC2), .y9(NET00004), .x10(WC_CSR0));
t398 cell_O24(.x1(WC_CSR0), .y2(NET00379), .x4(INIT3), .x5(nADC0), .x6(ADC0), .y9(NET00197), .x10(WC_CSR0));
t408 cell_M22(.q2(RD2), .q3(nRD2), .r5(NET00009), .s10(NET00011));
t376 cell_O21(.x1(nRP_DAT), .x3(nRD0), .y4(NET00129), .x6(nRC_DAT), .x8(nRD0), .y9(NET00371));
t376 cell_N8(.x1(nSA0), .x3(nDLA0), .y4(NET00370), .x6(SA1), .x8(HL0), .y9(NET00391));

endmodule
