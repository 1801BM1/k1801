//
// Copyright (c) 2013 by 1801BM1@gmail.com
//______________________________________________________________________________
//
`timescale 1ns / 100ps

module vp_120
(
   inout[9:0]  PIN_nADC,      // Central Address/Data inverted bus
                              //
   input       PIN_nSYNCC,    //
   input       PIN_nDINC,     //
   input       PIN_nDOUTC,    //
   input       PIN_nINITC,    //
   input       PIN_nCSC,      //
   output      PIN_nARC,      //
   output      PIN_nRPLYC,    //
                              //
   input       PIN_nIAKIC,    //
   output      PIN_nIAKOC,    //
   output      PIN_nVIRQC,    //
                              //
                              //
   inout[7:0]  PIN_nADP,      // Peripheral Address/Data inverted bus
                              //
   input       PIN_nSYNCP,    //
   input       PIN_nDINP,     //
   input       PIN_nDOUTP,    //
   input       PIN_nINITP,    //
   input       PIN_nCSP,      //
   output      PIN_nRPLYP,    //
                              //
   input       PIN_nIAKIP,    //
   output      PIN_nIAKOP,    //
   output      PIN_nVIRQP,    //
                              //
   output      PIN_A0,        //
   output      PIN_A1,        //
   output      PIN_nEP        //
);

//______________________________________________________________________________
//
// Autogenerated netlist
//
wire GND = 1'b0;
wire VCC = 1'b1;

wire nPT10;
wire CREQT1;
wire nPA04;
wire nCIET1;
wire CACKT1;
wire CACKT2;
wire nT11;
wire nT10;
wire PREQR1;
wire PACKRST;
wire PREQT0;
wire nPV7;
wire nT07;
wire INITC1;
wire CACKR1;
wire CACKR0;
wire nPR062;
wire nTRDY0;
wire nCW666;
wire TRDY1;
wire DOUTP;
wire PACKR0;
wire IRST;
wire nPIER0;
wire TRDY0M;
wire RRDY1;
wire nCIET0;
wire CACKT0;
wire PV2;
wire CREQR1;
wire nPW072;
wire nCA04;
wire nC177560;
wire nCR662;
wire nRRDY0;
wire nDINC;
wire DOUTC;
wire PDINOUT;
wire ADC6;
wire CA7;
wire nCA7;
wire nCA5;
wire nCA1;
wire CV4;
wire nADC6;
wire nCR660;
wire nCIER0;
wire nCIER1;
wire nC176670;
wire nCA9;
wire CV2;
wire INITC0;
wire nCA00;
wire nC176660;
wire nSYNCC0;
wire nSYNCP;
wire DINP;
wire nCSC;
wire nADP7;
wire nCSP;
wire PA1;
wire PMX0;
wire nT23;
wire PMX2;
wire nT22;
wire PMX1;
wire nPW070;
wire PA0;
wire nCR562;
wire CREQR0;
wire PREQRST;
wire nCA02;
wire PA2;
wire nPA00;
wire nPA2;
wire nPA06;
wire PA3;
wire nT00;
wire CA6;
wire nP177060;
wire nPA02;
wire nPA3;
wire PACKT1;
wire nPIER2;
wire PREQT1;
wire TRDY2;
wire CA2;
wire nCA6;
wire nADP2;
wire CREQT2;
wire CREQT0;
wire nADP6;
wire PACKR2;
wire nRRDY1;
wire nRSTIE;
wire PREQR2;
wire nDINP;
wire TRDY0;
wire nADP1;
wire CA9;
wire nCA4;
wire nPT12;
wire nPT11;
wire PACKT0;
wire nPIER1;
wire nPR064;
wire RRDY0;
wire nPR060;
wire nPR076;
wire nINITP;
wire DIS_CH0;
wire CA3;
wire nCA3;
wire nPT01;
wire nPT02;
wire PMX4;
wire PACKR1;
wire PV4;
wire nPIET1;
wire nCRSEL;
wire nT03;
wire CV8;
wire nCR560;
wire nCR664;
wire nCR674;
wire nTRDY1;
wire nPR066;
wire nP177070;
wire CSV7;
wire nCA06;
wire nCR564;
wire nT26;
wire nCW566;
wire nPIET0;
wire PV3;
wire PMX6;
wire PMX3;
wire PA6;
wire PA5;
wire PA4;
wire nPA1;
wire PA7;
wire nPA6;
wire nPA5;
wire INITP;
wire nPA4;
wire DINC;
wire nT25;
wire P177000;
wire C17XX60;
wire PV7;
wire PMX5;
wire nT24;
wire nPT13;
wire nPT14;
wire nT16;
wire nPT15;
wire nPT16;
wire nT15;
wire nT14;
wire nT06;
wire PV6;
wire nPT04;
wire nPT03;
wire PREQR0;
wire nPT05;
wire nT05;
wire CSV6;
wire nPT06;
wire CV5;
wire nT04;
wire nT13;
wire nCA2;
wire CA1;
wire nSYNCC;
wire nSYNCP0;
wire nCIET2;
wire nT02;
wire nT27;
wire nPT07;
wire nADP0;
wire ISET;
wire nPT17;
wire nPT00;
wire nT01;
wire nT12;
wire nT17;
wire nT20;
wire nT21;
wire PRPLY;
wire nCW676;
wire nTRDY2;

wire NET00000;
wire NET00001;
wire NET00002;
wire NET00004;
wire NET00006;
wire NET00009;
wire NET00012;
wire NET00013;
wire NET00014;
wire NET00016;
wire NET00018;
wire NET00019;
wire NET00020;
wire NET00021;
wire NET00024;
wire NET00026;
wire NET00029;
wire NET00030;
wire NET00033;
wire NET00032;
wire NET00039;
wire NET00040;
wire NET00041;
wire NET00042;
wire NET00047;
wire NET00050;
wire NET00051;
wire NET00052;
wire NET00053;
wire NET00056;
wire NET00207;
wire NET00060;
wire NET00065;
wire NET00066;
wire NET00067;
wire NET00068;
wire NET00069;
wire NET00071;
wire NET00073;
wire NET00075;
wire NET00080;
wire NET00083;
wire NET00084;
wire NET00089;
wire NET00092;
wire NET00096;
wire NET00097;
wire NET00098;
wire NET00100;
wire NET00104;
wire NET00105;
wire NET00110;
wire NET00111;
wire NET00112;
wire NET00117;
wire NET00118;
wire NET00120;
wire NET00122;
wire NET00123;
wire NET00124;
wire NET00125;
wire NET00506;
wire NET00128;
wire NET00130;
wire NET00131;
wire NET00132;
wire NET00133;
wire NET00134;
wire NET00136;
wire NET00138;
wire NET00139;
wire NET00140;
wire NET00142;
wire NET00144;
wire NET00510;
wire NET00146;
wire NET00151;
wire NET00152;
wire NET00153;
wire NET00154;
wire NET00160;
wire NET00166;
wire NET00168;
wire NET00513;
wire NET00172;
wire NET00514;
wire NET00175;
wire NET00176;
wire NET00177;
wire NET00178;
wire NET00198;
wire NET00226;
wire NET00184;
wire NET00185;
wire NET00188;
wire NET00189;
wire NET00192;
wire NET00196;
wire NET00227;
wire NET00256;
wire NET00199;
wire NET00201;
wire NET00203;
wire NET00204;
wire NET00206;
wire NET00264;
wire NET00208;
wire NET00210;
wire NET00211;
wire NET00212;
wire NET00216;
wire NET00217;
wire NET00218;
wire NET00219;
wire NET00286;
wire NET00221;
wire NET00222;
wire NET00295;
wire NET00224;
wire NET00225;
wire NET00296;
wire NET00360;
wire NET00228;
wire NET00361;
wire NET00232;
wire NET00234;
wire NET00362;
wire NET00239;
wire NET00386;
wire NET00242;
wire NET00387;
wire NET00245;
wire NET00248;
wire NET00390;
wire NET00252;
wire NET00254;
wire NET00255;
wire NET00393;
wire NET00257;
wire NET00261;
wire NET00263;
wire NET00265;
wire NET00266;
wire NET00268;
wire NET00269;
wire NET00270;
wire NET00271;
wire NET00272;
wire NET00412;
wire NET00275;
wire NET00276;
wire NET00277;
wire NET00414;
wire NET00282;
wire NET00283;
wire NET00285;
wire NET00415;
wire NET00287;
wire NET00288;
wire NET00289;
wire NET00291;
wire NET00418;
wire NET00297;
wire NET00299;
wire NET00300;
wire NET00301;
wire NET00302;
wire NET00303;
wire NET00305;
wire NET00420;
wire NET00307;
wire NET00421;
wire NET00313;
wire NET00316;
wire NET00317;
wire NET00318;
wire NET00422;
wire NET00327;
wire NET00425;
wire NET00330;
wire NET00334;
wire NET00335;
wire NET00336;
wire NET00337;
wire NET00426;
wire NET00339;
wire NET00340;
wire NET00427;
wire NET00342;
wire NET00343;
wire NET00344;
wire NET00346;
wire NET00347;
wire NET00348;
wire NET00349;
wire NET00353;
wire NET00354;
wire NET00435;
wire NET00359;
wire NET00363;
wire NET00447;
wire NET00366;
wire NET00367;
wire NET00368;
wire NET00371;
wire NET00372;
wire NET00448;
wire NET00449;
wire NET00379;
wire NET00380;
wire NET00381;
wire NET00383;
wire NET00384;
wire NET00399;
wire NET00400;
wire NET00401;
wire NET00402;
wire NET00411;
wire NET00481;
wire NET00398;
wire NET00483;
wire NET00484;
wire NET00485;
wire NET00486;
wire NET00487;
wire NET00405;
wire NET00406;
wire NET00488;
wire NET00489;
wire NET00490;
wire NET00495;
wire NET00497;
wire NET00413;
wire NET00501;
wire NET00515;
wire NET00516;
wire NET00471;
wire NET00474;
wire NET00475;
wire NET00477;
wire NET00431;
wire NET00432;
wire NET00467;
wire NET00478;
wire NET00436;
wire NET00465;
wire NET00464;
wire NET00498;
wire NET00458;
wire NET00511;
wire NET00507;
wire NET00457;
wire NET00456;
wire NET00517;
wire NET00502;
wire NET00500;

//______________________________________________________________________________
//
// Autogenerated cell instantiations
//
tOUTPUT_OE  cell_PINOU14(.x1(NET00218), .x2(NET00211), .y1(PIN_nADC[0]));
tOUTPUT_OE  cell_PINOU15(.x1(NET00219), .x2(NET00211), .y1(PIN_nADC[1]));
tOUTPUT_OE  cell_PINOU16(.x1(NET00221), .x2(NET00211), .y1(PIN_nADC[2]));
tOUTPUT_OE  cell_PINOU17(.x1(NET00222), .x2(NET00211), .y1(PIN_nADC[3]));
tOUTPUT_OE  cell_PINOU18(.x1(NET00210), .x2(NET00211), .y1(PIN_nADC[4]));
tOUTPUT_OE  cell_PINOU20(.x1(NET00349), .x2(NET00211), .y1(PIN_nADC[5]));
tOUTPUT_OE  cell_PINOU22(.x1(NET00348), .x2(NET00211), .y1(PIN_nADC[6]));
tOUTPUT_OE  cell_PINOU23(.x1(NET00347), .x2(NET00211), .y1(PIN_nADC[7]));
tOUTPUT_OE  cell_PINOU24(.x1(NET00346), .x2(NET00211), .y1(PIN_nADC[8]));

tINPUT      cell_PIN14(.y1(NET00144), .x1(PIN_nADC[0]));
tINPUT      cell_PIN15(.y1(NET00124), .x1(PIN_nADC[1]));
tINPUT      cell_PIN16(.y1(NET00245), .x1(PIN_nADC[2]));
tINPUT      cell_PIN17(.y1(NET00212), .x1(PIN_nADC[3]));
tINPUT      cell_PIN18(.y1(NET00178), .x1(PIN_nADC[4]));
tINPUT      cell_PIN20(.y1(NET00026), .x1(PIN_nADC[5]));
tINPUT      cell_PIN22(.y1(NET00020), .x1(PIN_nADC[6]));
tINPUT      cell_PIN23(.y1(NET00012), .x1(PIN_nADC[7]));
tINPUT      cell_PIN25(.y1(NET00208), .x1(PIN_nADC[9]));

tINPUT      cell_PIN9( .y2(NET00398), .x1(PIN_nINITC));
tINPUT      cell_PIN13(.y2(NET00405), .x1(PIN_nCSC));
tINPUT      cell_PIN6( .y1(nSYNCC0),  .x1(PIN_nSYNCC));
tINPUT      cell_PIN5( .y2(NET00112), .x1(PIN_nDINC));
tINPUT      cell_PIN4( .y2(NET00111), .x1(PIN_nDOUTC));
tINPUT      cell_PIN10(.y1(NET00068), .x1(PIN_nIAKIC));

tOUTPUT_OC  cell_PIN11(.x1(NET00406), .y1(PIN_nRPLYC));
tOUTPUT_OC  cell_PIN12(.x1(NET00380), .y1(PIN_nARC));
tOUTPUT_OC  cell_PIN19(.x1(NET00188), .y1(PIN_nVIRQC));
tOUTPUT     cell_PIN8( .x1(NET00498), .y1(PIN_nIAKOC));

tOUTPUT_OE  cell_PINOU3( .x1(NET00138), .x2(NET00030), .y1(PIN_nADP[0]));
tOUTPUT_OE  cell_PINOU2( .x1(NET00130), .x2(NET00030), .y1(PIN_nADP[1]));
tOUTPUT_OE  cell_PINOU1( .x1(NET00285), .x2(NET00030), .y1(PIN_nADP[2]));
tOUTPUT_OE  cell_PINOU40(.x1(NET00029), .x2(NET00030), .y1(PIN_nADP[3]));
tOUTPUT_OE  cell_PINOU39(.x1(NET00413), .x2(NET00030), .y1(PIN_nADP[4]));
tOUTPUT_OE  cell_PINOU38(.x1(NET00456), .x2(NET00030), .y1(PIN_nADP[5]));
tOUTPUT_OE  cell_PINOU37(.x1(NET00458), .x2(NET00030), .y1(PIN_nADP[6]));
tOUTPUT_OE  cell_PINOU36(.x1(NET00457), .x2(NET00030), .y1(PIN_nADP[7]));

tINPUT      cell_PIN3( .y1(nADP0),    .x1(PIN_nADP[0]));
tINPUT      cell_PIN2( .y1(nADP1),    .x1(PIN_nADP[1]));
tINPUT      cell_PIN1( .y1(nADP2),    .x1(PIN_nADP[2]));
tINPUT      cell_PIN40(.y1(NET00337), .x1(PIN_nADP[3]));
tINPUT      cell_PIN39(.y1(NET00128), .x1(PIN_nADP[4]));
tINPUT      cell_PIN38(.y1(NET00123), .x1(PIN_nADP[5]));
tINPUT      cell_PIN37(.y1(nADP6),    .x1(PIN_nADP[6]));
tINPUT      cell_PIN36(.y1(nADP7),    .x1(PIN_nADP[7]));

tINPUT      cell_PIN35(.y1(nINITP),   .x1(PIN_nINITP));
tINPUT      cell_PIN26(.y1(NET00297), .x1(PIN_nCSP));
tINPUT      cell_PIN30(.y1(nSYNCP0),  .x1(PIN_nSYNCP));
tINPUT      cell_PIN31(.y1(NET00092), .x1(PIN_nDINP));
tINPUT      cell_PIN32(.y1(NET00118), .x1(PIN_nDOUTP));
tINPUT      cell_PIN34(.y1(NET00047), .x1(PIN_nIAKIP));

tOUTPUT_OC  cell_PIN41(.x1(NET00500), .y1(PIN_nVIRQP));
tOUTPUT_OC  cell_PIN27(.x1(NET00291), .y1(PIN_nRPLYP));
tOUTPUT     cell_PIN7( .x1(NET00153), .y1(PIN_nIAKOP));

tOUTPUT     cell_PIN33(.x1(PA0),      .y1(PIN_A0));
tOUTPUT     cell_PIN28(.x1(PA1),      .y1(PIN_A1));
tOUTPUT     cell_PIN29(.x1(NET00305), .y1(PIN_nEP));

//______________________________________________________________________________
//
// t372 cell_A38(.x1(NET00475), .y2(NET00030), .y3(NET00030), .y4(NET00030), .x5(NET00475), .x6(NET00475));
t372 cell_A38(.x1(NET00475), .y2(NET00030), .x5(NET00475), .x6(NET00475));

t416 cell_A11(.c1(NET00160), .q3(CA2), .q4(nCA2), .d5(NET00245));
t376 cell_A1(.x1(CV5), .x3(NET00379), .y4(NET00381), .x6(NET00080), .x8(NET00380), .y9(NET00379));
t416 cell_A27(.c1(NET00248), .q4(nPT04), .d5(NET00128));
t416 cell_A19(.c1(NET00248), .q4(nPT01), .d5(nADP1));
t416 cell_A15(.c1(NET00248), .q4(nPT00), .d5(nADP0));
t390 cell_A3(.x1(CA1), .y4(nCA02), .x5(nCA2), .x6(nCA1), .y9(nCA00), .x10(nCA2));
t378 cell_A5(.x1(nCA5), .y2(NET00075), .x3(nCSC), .x5(nCA4));
t376 cell_A29(.x1(NET00110), .x3(nPT05), .y4(NET00383), .x6(NET00110), .x8(nPT04), .y9(NET00384));
t376 cell_A17(.x1(NET00110), .x3(nPT01), .y4(NET00252), .x6(NET00110), .x8(nPT00), .y9(NET00021));
t376 cell_A18(.x1(NET00217), .x3(NET00021), .y4(NET00218), .x6(NET00216), .x8(NET00252), .y9(NET00219));
t416 cell_A31(.c1(NET00248), .q4(nPT05), .d5(NET00123));
t416 cell_B19(.c1(NET00069), .q4(nPT11), .d5(nADP1));
t376 cell_A35(.x1(NET00110), .x3(nPT07), .y4(NET00471), .x6(NET00110), .x8(nPT06), .y9(NET00474));
t378 cell_A34(.x1(CSV6), .y2(NET00348), .x3(NET00465), .x5(NET00474));
t416 cell_B21(.c1(NET00069), .q4(nPT12), .d5(nADP2));
t380 cell_A36(.x1(CSV7), .y2(NET00346), .y3(NET00347), .x4(NET00464), .x5(CV8), .x6(NET00471));
t416 cell_A37(.c1(NET00248), .q4(nPT07), .d5(nADP7));
t376 cell_A23(.x1(NET00110), .x3(nPT03), .y4(NET00371), .x6(NET00110), .x8(nPT02), .y9(NET00372));
t378 cell_A24(.x1(CACKT2), .y2(NET00222), .x3(NET00353), .x5(NET00371));
t390 cell_A39(.x1(NET00477), .y4(NET00475), .x5(nPV7), .x6(P177000), .y9(NET00477), .x10(DINP));
t416 cell_A25(.c1(NET00248), .q4(nPT03), .d5(NET00337));
t416 cell_A21(.c1(NET00248), .q4(nPT02), .d5(nADP2));
t416 cell_A7(.c1(NET00160), .q3(CA1), .q4(nCA1), .d5(NET00124));
t376 cell_B17(.x1(NET00117), .x3(nPT11), .y4(NET00216), .x6(NET00117), .x8(nPT10), .y9(NET00217));
t416 cell_A33(.c1(NET00248), .q4(nPT06), .d5(nADP6));
t378 cell_A28(.x1(CV4), .y2(NET00210), .x3(NET00014), .x5(NET00384));
t378 cell_A30(.x1(CV5), .y2(NET00349), .x3(NET00359), .x5(NET00383));
t377 cell_B1(.x1(CV5), .y2(NET00380), .x3(NET00478), .y4(NET00406), .x5(NET00084), .x6(NET00083), .x8(NET00380), .y9(NET00478));
t378 cell_A22(.x1(CV2), .y2(NET00221), .x3(NET00354), .x5(NET00372));
t376 cell_B35(.x1(NET00117), .x3(nPT17), .y4(NET00464), .x6(NET00117), .x8(nPT16), .y9(NET00465));
t428 cell_E5(.x2(nSYNCC0), .y3(nSYNCC));
t374 cell_D1(.x1(C17XX60), .x2(nC176670), .x3(NET00263), .y4(nCRSEL), .y8(NET00263));
t381 cell_B5(.x1(CA9), .y2(NET00073), .x3(nCA7), .x4(nCA3), .x6(CA6));
t390 cell_B3(.x1(CA1), .y4(nCA06), .x5(CA2), .x6(nCA1), .y9(nCA04), .x10(CA2));
t390 cell_B39(.x1(P177000), .y4(NET00467), .x5(PDINOUT), .x6(NET00467), .y9(PRPLY), .x10(nPV7));
t416 cell_C19(.c1(NET00184), .q3(PA2), .q4(nPA2), .d5(nADP2));
t429 cell_E11(.y3(ADC6), .x5(NET00020));
t378 cell_D15(.x1(CREQR0), .y2(NET00154), .x3(CREQT0), .x5(CREQR1));
t379 cell_D9(.x1(CACKT2), .y2(NET00265), .x3(CACKT1), .y4(NET00266), .x5(CACKT0), .x6(CACKR0), .x8(CACKT0));
t429 cell_K0(.y3(nDINC), .x5(NET00112));
t416 cell_C31(.c1(NET00184), .q4(nCSP), .d5(NET00297));
t416 cell_C23(.c1(NET00184), .q3(PA4), .q4(nPA4), .d5(NET00128));
t428 cell_E25(.x2(NET00289), .y3(nP177070));
t390 cell_D17(.x1(PA1), .y4(nPA06), .x5(PA2), .x6(nPA1), .y9(nPA04), .x10(PA2));
t390 cell_D19(.x1(PA1), .y4(nPA02), .x5(nPA2), .x6(nPA1), .y9(nPA00), .x10(nPA2));
t428 cell_E1(.x2(NET00398), .y3(INITC1));
t416 cell_B25(.c1(NET00069), .q4(nPT13), .d5(NET00337));
t428 cell_E29(.x2(NET00303), .y3(nPR076));
t381 cell_D23(.x1(PA7), .y2(NET00316), .x3(PA6), .x4(nPA4), .x6(nPA5));
t390 cell_C3(.x1(NET00071), .y4(nC176660), .x5(NET00075), .x6(NET00073), .y9(nC176670), .x10(NET00075));
t391 cell_B9(.x1(NET00089), .x2(NET00265), .y3(CV2), .y4(CV5), .x5(NET00266), .x6(NET00089), .y9(CV4), .x10(NET00266));
t416 cell_C27(.c1(NET00184), .q3(PA6), .q4(nPA6), .d5(nADP6));
t429 cell_E33(.y3(DINP), .x5(NET00092));
t390 cell_D25(.x1(NET00316), .y4(NET00283), .x5(NET00317), .x6(NET00316), .y9(NET00289), .x10(NET00318));
t381 cell_D27(.x1(PA5), .y2(NET00313), .x3(PA4), .x4(PA2), .x6(PA3));
t416 cell_B13(.c1(NET00160), .q3(CA9), .q4(nCA9), .d5(NET00208));
t416 cell_B11(.c1(NET00160), .q3(CA3), .q4(nCA3), .d5(NET00212));
t376 cell_B29(.x1(NET00117), .x3(nPT15), .y4(NET00359), .x6(NET00117), .x8(nPT14), .y9(NET00014));
t428 cell_E37(.x2(nSYNCP0), .y3(nSYNCP));
t378 cell_D29(.x1(nCSP), .y2(NET00327), .x3(PA7), .x5(nPA6));
t416 cell_B15(.c1(NET00069), .q4(nPT10), .d5(nADP0));
t382 cell_G31(.x1(PACKR0), .y2(NET00363), .x3(PACKR1), .x4(PACKT0), .x5(NET00363), .x6(PACKT1), .y8(PV4));
t416 cell_B33(.c1(NET00069), .q4(nPT16), .d5(nADP6));
t388 cell_D31(.x1(NET00431), .y2(NET00431), .x3(NET00305), .y4(NET00432), .y5(NET00305), .x6(NET00313), .x7(PDINOUT), .x10(NET00327));
t378 cell_D33(.x1(nPA02), .y2(NET00232), .x3(nSYNCP), .x5(nP177060));
t374 cell_H37(.x1(NET00342), .x2(NET00343), .x3(NET00344), .y4(NET00343), .y8(PMX4));
t374 cell_I37(.x1(NET00334), .x2(NET00335), .x3(NET00336), .y4(NET00335), .y8(PMX1));
t376 cell_I39(.x1(DOUTP), .x3(DINP), .y4(NET00032), .x6(nSYNCP0), .x8(NET00032), .y9(PDINOUT));
t391 cell_H39(.x1(NET00339), .x2(NET00340), .y3(NET00242), .y4(NET00303), .x5(DINP), .x6(NET00339), .y9(NET00340), .x10(DOUTP));
t381 cell_C5(.x1(nCA7), .y2(NET00071), .x3(CA6), .x4(CA9), .x6(CA3));
t380 cell_C9(.x1(CACKT2), .y2(CV8), .y3(NET00089), .x4(CACKT1), .x5(NET00089), .x6(CACKR1));
t390 cell_D3(.x1(nC177560), .y4(C17XX60), .x5(nC176660), .x6(NET00261), .y9(nC177560), .x10(NET00075));
t416 cell_C13(.c1(NET00160), .q4(nCA4), .d5(NET00178));
t416 cell_D13(.c1(NET00160), .q3(CA6), .q4(nCA6), .d5(NET00020));
t378 cell_C35(.x1(nP177070), .y2(NET00302), .x3(nSYNCP), .x5(nPA00));
t378 cell_D35(.x1(nP177070), .y2(NET00234), .x3(nSYNCP), .x5(nPA02));
t389 cell_C37(.x1(nSYNCP), .x2(nPA00), .y3(NET00301), .x4(nP177060), .y5(P177000), .x6(nP177070), .x10(nP177060));
t378 cell_D37(.x1(nPA04), .y2(NET00201), .x3(nSYNCP), .x5(nP177060));
t378 cell_D39(.x1(nPA06), .y2(NET00366), .x3(nSYNCP), .x5(nP177060));
t373 cell_J37(.x1(nPR066), .x3(nPIER2), .y4(PMX2));
t381 cell_H31(.x1(PACKRST), .y2(NET00330), .x3(PACKR0), .x4(PACKR1), .x6(PACKR2));
t390 cell_J39(.x1(NET00301), .y4(nPR060), .x5(DINP), .x6(DOUTP), .y9(nPW070), .x10(NET00302));
t378 cell_H29(.x1(nDINP), .y2(PACKT1), .x3(NET00192), .x5(NET00177));
t390 cell_L39(.x1(NET00232), .y4(nPR062), .x5(DINP), .x6(NET00234), .y9(nPW072), .x10(DOUTP));
t377 cell_C1(.x1(DINC), .y2(NET00080), .x3(DOUTC), .y4(NET00083), .x5(DINC), .x6(nCRSEL), .x8(nSYNCC0), .y9(NET00084));
t416 cell_B7(.c1(NET00160), .q3(nCSC), .d5(NET00405));
t428 cell_E0(.x2(NET00398), .y3(INITC0));
t416 cell_B37(.c1(NET00069), .q4(nPT17), .d5(nADP7));
t416 cell_C33(.c1(NET00184), .q3(PA0), .d5(nADP0));
t416 cell_C29(.c1(NET00184), .q3(PA7), .d5(nADP7));
t416 cell_C17(.c1(NET00184), .q3(PA1), .q4(nPA1), .d5(nADP1));
t376 cell_B23(.x1(NET00117), .x3(nPT13), .y4(NET00353), .x6(NET00117), .x8(nPT12), .y9(NET00354));
t416 cell_C21(.c1(NET00184), .q3(PA3), .q4(nPA3), .d5(NET00337));
t416 cell_C25(.c1(NET00184), .q3(PA5), .q4(nPA5), .d5(NET00123));
t428 cell_E7(.x2(NET00381), .y3(NET00211));
t428 cell_E27(.x2(NET00283), .y3(nP177060));
t429 cell_E13(.y3(nADC6), .x5(ADC6));
t428 cell_E31(.x2(NET00368), .y3(nPR066));
t376 cell_D21(.x1(PA3), .x3(nCSP), .y4(NET00317), .x6(nCSP), .x8(nPA3), .y9(NET00318));
t406 cell_F21(.c1(VCC), .r2(INITC0), .q3(NET00257), .r5(RRDY0), .s10(PACKT0));
t378 cell_F1(.x1(nC177560), .y2(NET00483), .x3(nSYNCC), .x5(nCA00));
t389 cell_H8(.x1(NET00268), .x2(NET00270), .y3(NET00269), .x4(NET00272), .y5(CSV7), .x6(NET00269), .x10(NET00271));
t416 cell_G13(.c1(nDINC), .q3(NET00039), .q4(NET00040), .d5(CREQT0));
t391 cell_H3(.x1(NET00275), .x2(NET00277), .y3(NET00276), .y4(NET00277), .x5(DOUTC), .x6(DINC), .y9(nCR660), .x10(NET00275));
t376 cell_J7(.x1(NET00282), .x3(NET00490), .y4(NET00271), .x6(nCR674), .x8(TRDY2), .y9(NET00490));
t391 cell_F3(.x1(NET00483), .x2(NET00484), .y3(NET00481), .y4(NET00484), .x5(DOUTC), .x6(DINC), .y9(nCR560), .x10(NET00483));
t406 cell_F5(.c1(NET00481), .r2(INITC1), .q4(nCIER0), .r5(nADC6), .s10(ADC6));
t378 cell_I9(.x1(nDINC), .y2(CACKT1), .x3(NET00399), .x5(NET00002));
t416 cell_I13(.c1(nDINC), .q3(NET00399), .q4(NET00516), .d5(CREQT1));
t391 cell_J3(.x1(NET00487), .x2(NET00489), .y3(NET00488), .y4(NET00489), .x5(DOUTC), .x6(DINC), .y9(nCR674), .x10(NET00487));
t378 cell_G1(.x1(nC177560), .y2(NET00104), .x3(nSYNCC), .x5(nCA04));
t378 cell_J9(.x1(nDINC), .y2(CACKT2), .x3(NET00486), .x5(NET00485));
t374 cell_G6(.x1(TRDY0), .x2(NET00098), .x3(nCIET0), .y4(NET00098), .y8(TRDY0M));
t428 cell_K3(.x2(NET00111), .y3(DOUTC));
t378 cell_L3(.x1(nCA06), .y2(NET00300), .x3(nC177560), .x5(nSYNCC));
t378 cell_I1(.x1(nC176660), .y2(NET00400), .x3(nSYNCC), .x5(nCA04));
t406 cell_I5(.c1(NET00401), .r2(INITC1), .q4(nCIET1), .r5(nADC6), .s10(ADC6));
t428 cell_K9(.x2(nCR662), .y3(NET00110));
t428 cell_K5(.x2(nCR562), .y3(NET00117));
t384 cell_O3(.x1(NET00146), .y3(nCW676), .x5(DOUTC));
t376 cell_F7(.x1(nCR560), .x3(nRRDY0), .y4(NET00270), .x6(nCR564), .x8(TRDY0), .y9(NET00272));
t378 cell_M1(.x1(nCA02), .y2(NET00411), .x3(nC176660), .x5(nSYNCC));
t378 cell_L1(.x1(nCA02), .y2(NET00299), .x3(nC177560), .x5(nSYNCC));
t429 cell_K11(.y3(NET00436), .x5(nCW666));
t390 cell_N3(.x1(NET00501), .y4(nCW666), .x5(DOUTC), .x6(NET00411), .y9(nCR662), .x10(DINC));
t376 cell_H7(.x1(nCR660), .x3(nRRDY1), .y4(NET00282), .x6(nCR664), .x8(TRDY1), .y9(NET00268));
t378 cell_N1(.x1(nCA06), .y2(NET00501), .x3(nC176660), .x5(nSYNCC));
t378 cell_O1(.x1(nC176670), .y2(NET00146), .x3(nSYNCC), .x5(nCA06));
t378 cell_F9(.x1(nDINC), .y2(CACKR0), .x3(NET00065), .x5(NET00068));
t380 cell_G11(.x1(NET00042), .y2(NET00001), .y3(NET00041), .x4(NET00040), .x5(NET00041), .x6(nDINC));
t380 cell_H11(.x1(NET00001), .y2(NET00002), .y3(NET00000), .x4(NET00004), .x5(NET00000), .x6(nDINC));
t378 cell_F15(.x1(nCIER0), .y2(CREQR0), .x3(NET00060), .x5(nRRDY0));
t378 cell_G9(.x1(nDINC), .y2(CACKT0), .x3(NET00039), .x5(NET00042));
t391 cell_G3(.x1(DOUTC), .x2(NET00105), .y3(NET00100), .y4(NET00105), .x5(NET00104), .x6(DINC), .y9(nCR564), .x10(NET00104));
t378 cell_H9(.x1(nDINC), .y2(CACKR1), .x3(NET00006), .x5(NET00001));
t380 cell_I11(.x1(NET00002), .y2(NET00485), .y3(NET00515), .x4(NET00516), .x5(NET00515), .x6(nDINC));
t416 cell_F13(.c1(nDINC), .q3(NET00065), .q4(NET00066), .d5(CREQR0));
t376 cell_I7(.x1(nCR660), .x3(nCIER1), .y4(NET00287), .x6(nCR664), .x8(nCIET1), .y9(NET00288));
t378 cell_H1(.x1(nC176660), .y2(NET00275), .x3(nSYNCC), .x5(nCA00));
t378 cell_J1(.x1(nC176670), .y2(NET00487), .x3(nSYNCC), .x5(nCA04));
t406 cell_G5(.c1(NET00100), .r2(INITC1), .q4(nCIET0), .r5(nADC6), .s10(ADC6));
t406 cell_H5(.c1(NET00276), .r2(INITC1), .q4(nCIER1), .r5(nADC6), .s10(ADC6));
t406 cell_J5(.c1(NET00488), .r2(INITC1), .q4(nCIET2), .r5(nADC6), .s10(ADC6));
t429 cell_K7(.y3(NET00013), .x5(nCW566));
t380 cell_J11(.x1(NET00485), .y2(NET00498), .y3(NET00497), .x4(NET00495), .x5(NET00497), .x6(nDINC));
t416 cell_H13(.c1(nDINC), .q3(NET00006), .q4(NET00004), .d5(CREQR1));
t391 cell_I3(.x1(NET00400), .x2(NET00402), .y3(NET00401), .y4(NET00402), .x5(DOUTC), .x6(DINC), .y9(nCR664), .x10(NET00400));
t416 cell_J13(.c1(nDINC), .q3(NET00486), .q4(NET00495), .d5(CREQT2));
t390 cell_M3(.x1(NET00300), .y4(nCW566), .x5(DOUTC), .x6(NET00299), .y9(nCR562), .x10(DINC));
t428 cell_K1(.x2(NET00112), .y3(DINC));
t376 cell_G7(.x1(nCR560), .x3(nCIER0), .y4(NET00096), .x6(nCR564), .x8(nCIET0), .y9(NET00097));
t429 cell_K13(.y3(NET00125), .x5(nCW676));
t380 cell_F11(.x1(NET00068), .y2(NET00042), .y3(NET00067), .x4(NET00066), .x5(NET00067), .x6(nDINC));
t411 cell_F19(.q1(RRDY0), .r3(INITC0), .q4(nRRDY0), .r5(nCR562), .s10(nPW070));
t381 cell_L9(.x1(NET00097), .y2(NET00286), .x3(NET00287), .x4(NET00096), .x6(NET00288));
t411 cell_G19(.q1(TRDY0), .r3(INITC0), .q4(nTRDY0), .r5(nPR060), .s10(nCW566));
t411 cell_H19(.q1(RRDY1), .r3(INITC0), .q4(nRRDY1), .r5(nCR662), .s10(nPW072));
t416 cell_M9(.c1(NET00013), .q4(nT01), .d5(NET00124));
t416 cell_N9(.c1(NET00436), .q4(nT11), .d5(NET00124));
t411 cell_I19(.q1(TRDY1), .r3(INITC0), .q4(nTRDY1), .r5(nPR062), .s10(nCW666));
t402 cell_G21(.r1(nTRDY0), .q3(NET00228), .s6(PACKR0));
t378 cell_F23(.x1(nPIET0), .y2(PREQT0), .x3(NET00257), .x5(RRDY0));
t378 cell_G23(.x1(nPIER0), .y2(PREQR0), .x3(NET00228), .x5(nTRDY0));
t380 cell_J27(.x1(NET00120), .y2(NET00153), .y3(NET00152), .x4(NET00151), .x5(NET00152), .x6(nDINP));
t406 cell_H21(.c1(VCC), .r2(INITC0), .q3(NET00196), .r5(RRDY1), .s10(PACKT1));
t416 cell_F25(.c1(nDINP), .q3(NET00254), .q4(NET00255), .d5(PREQT0));
t416 cell_H25(.c1(nDINP), .q3(NET00192), .q4(NET00199), .d5(PREQT1));
t416 cell_G25(.c1(nDINP), .q3(NET00224), .q4(NET00225), .d5(PREQR0));
t411 cell_J19(.q1(TRDY2), .r3(INITC0), .q4(nTRDY2), .r5(nPR064), .s10(nCW676));
t416 cell_M11(.c1(NET00013), .q4(nT02), .d5(NET00245));
t416 cell_O9(.c1(NET00125), .q4(nT21), .d5(NET00124));
t378 cell_F29(.x1(nDINP), .y2(PACKT0), .x3(NET00254), .x5(NET00227));
t380 cell_F31(.x1(PACKT1), .y2(PV3), .y3(NET00393), .x4(PACKR1), .x5(NET00393), .x6(PACKRST));
t416 cell_N11(.c1(NET00436), .q4(nT12), .d5(NET00245));
t402 cell_I21(.r1(nTRDY1), .q3(NET00172), .s6(PACKR1));
t378 cell_I23(.x1(nPIER1), .y2(PREQR1), .x3(NET00172), .x5(nTRDY1));
t378 cell_H23(.x1(nPIET1), .y2(PREQT1), .x3(NET00196), .x5(RRDY1));
t378 cell_J23(.x1(nPIER2), .y2(PREQR2), .x3(NET00142), .x5(nTRDY2));
t402 cell_J21(.r1(nTRDY2), .q3(NET00142), .s6(PACKR2));
t402 cell_H17(.r1(nRRDY1), .q3(NET00009), .s6(CACKR1));
t416 cell_O11(.c1(NET00125), .q4(nT22), .d5(NET00245));
t376 cell_F35(.x1(nPR076), .x3(RRDY0), .y4(NET00386), .x6(nPR066), .x8(nTRDY0), .y9(NET00387));
t406 cell_F33(.c1(NET00242), .r2(INITP), .q4(nPIET0), .r5(nADP0), .s10(NET00206));
t383 cell_O14(.x1(PV3), .y2(NET00029), .x3(NET00420), .x4(NET00422), .x5(PMX3), .x6(NET00421));
t383 cell_O12(.x1(PV2), .y2(NET00285), .x3(NET00425), .x4(NET00427), .x5(PMX2), .x6(NET00426));
t378 cell_F39(.x1(nP177070), .y2(NET00339), .x3(nSYNCP), .x5(nPA06));
t383 cell_D5(.x1(nCA9), .y2(NET00261), .x3(CA7), .x4(nCA6), .x5(DIS_CH0), .x6(CA3));
t391 cell_G39(.x1(NET00366), .x2(NET00367), .y3(NET00239), .y4(NET00368), .x5(DINP), .x6(NET00366), .y9(NET00367), .x10(DOUTP));
t416 cell_B31(.c1(NET00069), .q4(nPT15), .d5(NET00123));
t416 cell_B27(.c1(NET00069), .q4(nPT14), .d5(NET00128));
t428 cell_E39(.x2(nSYNCP0), .y3(NET00184));
t378 cell_J29(.x1(nDINP), .y2(PACKR2), .x3(NET00122), .x5(NET00120));
t384 cell_M39(.x1(NET00201), .y3(nPR064), .x5(DINP));
t416 cell_M5(.c1(NET00013), .q4(nT00), .d5(NET00144));
t374 cell_F37(.x1(NET00387), .x2(NET00390), .x3(NET00386), .y4(NET00390), .y8(PMX3));
t376 cell_N13(.x1(NET00264), .x3(nT13), .y4(NET00422), .x6(NET00264), .x8(nT12), .y9(NET00427));
t376 cell_O13(.x1(NET00134), .x3(nT23), .y4(NET00421), .x6(NET00134), .x8(nT22), .y9(NET00426));
t376 cell_M27(.x1(NET00016), .x3(nT07), .y4(NET00018), .x6(NET00016), .x8(nT06), .y9(NET00019));
t429 cell_K33(.y3(INITP), .x5(nINITP));
t381 cell_O8(.x1(PMX1), .y2(NET00130), .x3(NET00131), .x4(NET00133), .x6(NET00132));
t429 cell_E35(.y3(DOUTP), .x5(NET00118));
t428 cell_E3(.x2(nSYNCC0), .y3(NET00160));
t391 cell_I31(.x1(NET00307), .x2(PV7), .y3(nPV7), .y4(PV7), .x5(NET00330), .x6(NET00330), .y9(PV6), .x10(NET00307));
t416 cell_C11(.c1(NET00160), .q4(nCA5), .d5(NET00026));
t416 cell_D11(.c1(NET00160), .q3(CA7), .q4(nCA7), .d5(NET00012));
t406 cell_H33(.c1(NET00242), .r2(INITP), .q4(nPIET1), .r5(nADP1), .s10(NET00204));
t416 cell_O5(.c1(NET00125), .q4(nT20), .d5(NET00144));
t380 cell_J31(.x1(PACKT1), .y2(PV2), .y3(NET00307), .x4(PACKT0), .x5(NET00307), .x6(INITP));
t381 cell_O6(.x1(PMX0), .y2(NET00138), .x3(NET00139), .x4(NET00140), .x6(NET00136));
t416 cell_M15(.c1(NET00013), .q4(nT03), .d5(NET00212));
t376 cell_N27(.x1(NET00264), .x3(nT17), .y4(NET00507), .x6(NET00264), .x8(nT16), .y9(NET00511));
t429 cell_K37(.y3(NET00248), .x5(nPW072));
t376 cell_M7(.x1(NET00016), .x3(nT01), .y4(NET00131), .x6(NET00016), .x8(nT00), .y9(NET00139));
t388 cell_C15(.x1(CREQT1), .y2(NET00188), .x3(CREQT2), .y4(NET00189), .y5(NET00185), .x6(NET00154), .x7(NET00185), .x10(NET00189));
t373 cell_C39(.x1(NET00432), .x3(PRPLY), .y4(NET00291));
t373 cell_J35(.x1(nPR066), .x3(nTRDY2), .y4(PMX5));
t378 cell_G29(.x1(nDINP), .y2(PACKR0), .x3(NET00224), .x5(NET00052));
t378 cell_I29(.x1(nDINP), .y2(PACKR1), .x3(NET00168), .x5(NET00166));
t428 cell_K27(.x2(NET00092), .y3(nDINP));
t428 cell_K31(.x2(nPR060), .y3(NET00016));
t406 cell_G33(.c1(NET00239), .r2(INITP), .q4(nPIER0), .r5(nADP0), .s10(NET00206));
t416 cell_N5(.c1(NET00436), .q4(nT10), .d5(NET00144));
t388 cell_L7(.x1(nCIET2), .y2(NET00295), .x3(nCR674), .y4(NET00296), .y5(CSV6), .x6(NET00286), .x7(NET00296), .x10(NET00295));
t376 cell_O7(.x1(NET00134), .x3(nT21), .y4(NET00132), .x6(NET00134), .x8(nT20), .y9(NET00136));
t416 cell_I25(.c1(nDINP), .q3(NET00168), .q4(NET00176), .d5(PREQR1));
t406 cell_F17(.c1(VCC), .r2(nCIER0), .q3(NET00060), .r5(nRRDY0), .s10(CACKR0));
t416 cell_N15(.c1(NET00436), .q4(nT13), .d5(NET00212));
t380 cell_F27(.x1(NET00227), .y2(NET00166), .y3(NET00256), .x4(NET00255), .x5(NET00256), .x6(nDINP));
t406 cell_G17(.c1(VCC), .r2(TRDY0M), .q3(NET00033), .r5(INITC0), .s10(CACKT0));
t378 cell_H15(.x1(nCIER1), .y2(CREQR1), .x3(NET00009), .x5(nRRDY1));
t416 cell_M17(.c1(NET00013), .q4(nT04), .d5(NET00178));
t380 cell_H27(.x1(NET00177), .y2(NET00120), .y3(NET00198), .x4(NET00199), .x5(NET00198), .x6(nDINP));
t380 cell_I27(.x1(NET00176), .y2(NET00177), .y3(NET00175), .x4(NET00166), .x5(NET00175), .x6(nDINP));
t378 cell_I15(.x1(nCIET1), .y2(CREQT1), .x3(NET00517), .x5(TRDY1));
t378 cell_J15(.x1(nCIET2), .y2(CREQT2), .x3(NET00502), .x5(TRDY2));
t416 cell_N17(.c1(NET00436), .q4(nT14), .d5(NET00178));
t406 cell_I33(.c1(NET00239), .r2(INITP), .q4(nPIER1), .r5(nADP1), .s10(NET00204));
t406 cell_J33(.c1(NET00239), .r2(INITP), .q4(nPIER2), .r5(nADP2), .s10(NET00203));
t383 cell_O18(.x1(PV4), .y2(NET00413), .x3(NET00412), .x4(NET00415), .x5(PMX4), .x6(NET00414));
t376 cell_G35(.x1(nPR076), .x3(nPIET0), .y4(NET00360), .x6(nPR066), .x8(nPIER0), .y9(NET00361));
t376 cell_H35(.x1(nPR076), .x3(RRDY1), .y4(NET00344), .x6(nPR066), .x8(nTRDY1), .y9(NET00342));
t402 cell_M19(.r1(NET00448), .q3(NET00449), .s6(IRST));
t376 cell_N19(.x1(NET00264), .x3(nT15), .y4(NET00435), .x6(NET00264), .x8(nT14), .y9(NET00415));
t374 cell_G37(.x1(NET00361), .x2(NET00362), .x3(NET00360), .y4(NET00362), .y8(PMX0));
t376 cell_O19(.x1(NET00134), .x3(nT25), .y4(NET00418), .x6(NET00134), .x8(nT24), .y9(NET00414));
t383 cell_O20(.x1(PACKR2), .y2(NET00456), .x3(NET00447), .x4(NET00435), .x5(PMX5), .x6(NET00418));
t416 cell_M21(.c1(NET00013), .q4(nT05), .d5(NET00026));
t428 cell_K39(.x2(nPR064), .y3(NET00134));
t428 cell_K35(.x2(nPR062), .y3(NET00264));
t429 cell_K29(.y3(NET00069), .x5(nPW070));
t376 cell_N7(.x1(NET00264), .x3(nT11), .y4(NET00133), .x6(NET00264), .x8(nT10), .y9(NET00140));
t376 cell_M13(.x1(NET00016), .x3(nT03), .y4(NET00420), .x6(NET00016), .x8(nT02), .y9(NET00425));
t380 cell_L27(.x1(NET00047), .y2(NET00052), .y3(NET00051), .x4(NET00053), .x5(NET00051), .x6(nDINP));
t416 cell_J25(.c1(nDINP), .q3(NET00122), .q4(NET00151), .d5(PREQR2));
t380 cell_G27(.x1(NET00052), .y2(NET00227), .y3(NET00226), .x4(NET00225), .x5(NET00226), .x6(nDINP));
t416 cell_N21(.c1(NET00436), .q4(nT15), .d5(NET00026));
t378 cell_L23(.x1(nRSTIE), .y2(PREQRST), .x3(NET00056), .x5(ISET));
t378 cell_N23(.x1(PREQR1), .y2(NET00513), .x3(PREQT1), .x5(PREQR2));
t385 cell_O23(.x1(NET00513), .x2(NET00514), .y3(NET00514), .x5(NET00024), .y8(NET00500));
t416 cell_M25(.c1(NET00013), .q4(nT06), .d5(NET00020));
t416 cell_L25(.c1(nDINP), .q3(NET00050), .q4(NET00053), .d5(PREQRST));
t416 cell_N25(.c1(NET00436), .q4(nT16), .d5(NET00020));
t416 cell_O25(.c1(NET00125), .q4(nT26), .d5(NET00020));
t383 cell_O26(.x1(PV6), .y2(NET00458), .x3(NET00019), .x4(NET00511), .x5(PMX6), .x6(NET00510));
t376 cell_O27(.x1(NET00134), .x3(nT27), .y4(NET00506), .x6(NET00134), .x8(nT26), .y9(NET00510));
t378 cell_L29(.x1(nDINP), .y2(PACKRST), .x3(NET00050), .x5(NET00047));
t376 cell_M18(.x1(NET00016), .x3(nT05), .y4(NET00447), .x6(NET00016), .x8(nT04), .y9(NET00412));
t416 cell_O17(.c1(NET00125), .q4(nT24), .d5(NET00178));
t416 cell_O15(.c1(NET00125), .q4(nT23), .d5(NET00212));
t416 cell_M29(.c1(NET00013), .q4(nT07), .d5(NET00012));
t416 cell_O29(.c1(NET00125), .q4(nT27), .d5(NET00012));
t371 cell_M33(.x1(nADP0), .y3(NET00206), .y4(NET00207), .x6(nADP6));
t373 cell_L35(.x1(nRSTIE), .x3(nPR066), .y4(PMX6));
t371 cell_M35(.x1(nADP2), .y3(NET00203), .y4(NET00204), .x6(nADP1));
t416 cell_O21(.c1(NET00125), .q4(nT25), .d5(NET00026));
t378 cell_M23(.x1(PREQRST), .y2(NET00024), .x3(PREQR0), .x5(PREQT0));
t381 cell_O28(.x1(PV7), .y2(NET00457), .x3(NET00018), .x4(NET00507), .x6(NET00506));
t416 cell_N29(.c1(NET00436), .q4(nT17), .d5(NET00012));
t406 cell_L33(.c1(NET00239), .r2(INITP), .q4(nRSTIE), .r5(nADP6), .s10(NET00207));
t406 cell_L31(.c1(NET00242), .r2(INITP), .q3(DIS_CH0), .r5(nADP2), .s10(NET00203));
t378 cell_G15(.x1(GND), .y2(CREQT0), .x3(NET00033), .x5(TRDY0M));
t377 cell_L19(.x1(nINITP), .y2(NET00448), .x3(NET00448), .y4(IRST), .x5(INITC0), .x6(NET00448), .x8(NET00449), .y9(ISET));
t376 cell_I35(.x1(nPR076), .x3(nPIET1), .y4(NET00336), .x6(nPR066), .x8(nPIER1), .y9(NET00334));
t406 cell_L21(.c1(VCC), .r2(IRST), .q4(NET00056), .r5(PACKRST), .s10(ISET));
t406 cell_I17(.c1(VCC), .r2(TRDY1), .q3(NET00517), .r5(INITC0), .s10(CACKT1));
t406 cell_J17(.c1(VCC), .r2(TRDY2), .q3(NET00502), .r5(INITC0), .s10(CACKT2));
endmodule
